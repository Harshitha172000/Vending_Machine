VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vm
  CLASS BLOCK ;
  FOREIGN vm ;
  ORIGIN 0.000 0.000 ;
  SIZE 112.945 BY 123.665 ;
  PIN change[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END change[0]
  PIN change[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 119.665 109.850 123.665 ;
    END
  END change[1]
  PIN choice[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END choice[0]
  PIN choice[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END choice[1]
  PIN choice[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.945 73.480 112.945 74.080 ;
    END
  END choice[2]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 119.665 16.930 123.665 ;
    END
  END clk
  PIN coin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END coin[0]
  PIN coin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END coin[1]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.945 27.240 112.945 27.840 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 119.665 79.490 123.665 ;
    END
  END out[2]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 119.665 48.210 123.665 ;
    END
  END reset
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 89.435 10.640 91.035 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 55.550 10.640 57.150 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.665 10.640 23.265 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 93.705 107.180 95.305 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 60.160 107.180 61.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.615 107.180 28.215 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 72.495 10.640 74.095 111.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 38.605 10.640 40.205 111.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 76.935 107.180 78.535 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 43.385 107.180 44.985 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 107.180 111.605 ;
      LAYER met1 ;
        RECT 2.830 10.640 109.870 111.760 ;
      LAYER met2 ;
        RECT 2.860 119.385 16.370 119.665 ;
        RECT 17.210 119.385 47.650 119.665 ;
        RECT 48.490 119.385 78.930 119.665 ;
        RECT 79.770 119.385 109.290 119.665 ;
        RECT 2.860 4.280 109.840 119.385 ;
        RECT 3.410 4.000 32.930 4.280 ;
        RECT 33.770 4.000 64.210 4.280 ;
        RECT 65.050 4.000 95.490 4.280 ;
        RECT 96.330 4.000 109.840 4.280 ;
      LAYER met3 ;
        RECT 4.000 96.240 108.945 111.685 ;
        RECT 4.400 94.840 108.945 96.240 ;
        RECT 4.000 74.480 108.945 94.840 ;
        RECT 4.000 73.080 108.545 74.480 ;
        RECT 4.000 50.000 108.945 73.080 ;
        RECT 4.400 48.600 108.945 50.000 ;
        RECT 4.000 28.240 108.945 48.600 ;
        RECT 4.000 26.840 108.545 28.240 ;
        RECT 4.000 10.715 108.945 26.840 ;
      LAYER met4 ;
        RECT 23.665 10.640 38.205 111.760 ;
        RECT 40.605 10.640 55.150 111.760 ;
        RECT 57.550 10.640 72.095 111.760 ;
      LAYER met5 ;
        RECT 5.520 63.360 107.180 75.335 ;
        RECT 5.520 46.585 107.180 58.560 ;
        RECT 5.520 29.815 107.180 41.785 ;
  END
END vm
END LIBRARY

