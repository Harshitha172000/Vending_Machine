magic
tech sky130A
magscale 1 2
timestamp 1619947779
<< obsli1 >>
rect 1104 2159 11960 13073
<< obsm1 >>
rect 1104 1912 11960 13104
<< metal2 >>
rect 3238 0 3294 200
rect 9770 0 9826 200
<< obsm2 >>
rect 1398 256 11022 13705
rect 1398 200 3182 256
rect 3350 200 9714 256
rect 9882 200 11022 256
<< metal3 >>
rect 0 13608 200 13728
rect 12902 13608 13102 13728
rect 0 10616 200 10736
rect 12902 10616 13102 10736
rect 0 7488 200 7608
rect 12902 7488 13102 7608
rect 0 4496 200 4616
rect 12902 4496 13102 4616
rect 0 1504 200 1624
rect 12902 1504 13102 1624
<< obsm3 >>
rect 280 13528 12822 13701
rect 200 10816 12902 13528
rect 280 10536 12822 10816
rect 200 7688 12902 10536
rect 280 7408 12822 7688
rect 200 4696 12902 7408
rect 280 4416 12822 4696
rect 200 1704 12902 4416
rect 280 1531 12822 1704
<< metal4 >>
rect 2753 2128 3073 13104
rect 4563 2128 4883 13104
rect 6372 2128 6692 13104
rect 8181 2128 8501 13104
rect 9991 2128 10311 13104
<< obsm4 >>
rect 4107 2128 4483 13104
rect 4963 2128 6292 13104
rect 6772 2128 8101 13104
rect 8581 2128 9911 13104
<< metal5 >>
rect 1104 11035 11960 11355
rect 1104 9221 11960 9541
rect 1104 7408 11960 7728
rect 1104 5595 11960 5915
rect 1104 3781 11960 4101
<< obsm5 >>
rect 1104 9861 11960 10715
rect 1104 8048 11960 8901
rect 1104 6235 11960 7088
<< labels >>
rlabel metal3 s 12902 10616 13102 10736 6 change[0]
port 1 nsew signal output
rlabel metal3 s 12902 13608 13102 13728 6 change[1]
port 2 nsew signal output
rlabel metal3 s 0 1504 200 1624 6 choice[0]
port 3 nsew signal input
rlabel metal3 s 0 4496 200 4616 6 choice[1]
port 4 nsew signal input
rlabel metal3 s 0 7488 200 7608 6 choice[2]
port 5 nsew signal input
rlabel metal2 s 3238 0 3294 200 6 clk
port 6 nsew signal input
rlabel metal3 s 0 10616 200 10736 6 coin[0]
port 7 nsew signal input
rlabel metal3 s 0 13608 200 13728 6 coin[1]
port 8 nsew signal input
rlabel metal3 s 12902 1504 13102 1624 6 out[0]
port 9 nsew signal output
rlabel metal3 s 12902 4496 13102 4616 6 out[1]
port 10 nsew signal output
rlabel metal3 s 12902 7488 13102 7608 6 out[2]
port 11 nsew signal output
rlabel metal2 s 9770 0 9826 200 6 reset
port 12 nsew signal input
rlabel metal4 s 9991 2128 10311 13104 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 13104 6 VPWR
port 14 nsew power bidirectional
rlabel metal4 s 2753 2128 3073 13104 6 VPWR
port 15 nsew power bidirectional
rlabel metal5 s 1104 11035 11960 11355 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1104 7408 11960 7728 6 VPWR
port 17 nsew power bidirectional
rlabel metal5 s 1104 3781 11960 4101 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 8181 2128 8501 13104 6 VGND
port 19 nsew ground bidirectional
rlabel metal4 s 4563 2128 4883 13104 6 VGND
port 20 nsew ground bidirectional
rlabel metal5 s 1104 9221 11960 9541 6 VGND
port 21 nsew ground bidirectional
rlabel metal5 s 1104 5595 11960 5915 6 VGND
port 22 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 13102 13728
string LEFview TRUE
<< end >>
