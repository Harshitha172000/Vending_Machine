magic
tech sky130A
magscale 1 2
timestamp 1619947793
<< checkpaint >>
rect -3932 -3932 17034 17660
<< locali >>
rect 8493 9911 8527 10149
rect 6561 9503 6595 9673
rect 3617 8483 3651 8585
rect 7389 7395 7423 7497
<< viali >>
rect 4169 12801 4203 12835
rect 4077 12733 4111 12767
rect 4353 12733 4387 12767
rect 4813 12665 4847 12699
rect 2237 12257 2271 12291
rect 2329 12257 2363 12291
rect 5733 12257 5767 12291
rect 7665 12257 7699 12291
rect 8217 12257 8251 12291
rect 4905 12189 4939 12223
rect 5457 12189 5491 12223
rect 5917 12189 5951 12223
rect 8677 12189 8711 12223
rect 7757 12121 7791 12155
rect 2053 12053 2087 12087
rect 2513 12053 2547 12087
rect 3433 11849 3467 11883
rect 9965 11781 9999 11815
rect 4445 11713 4479 11747
rect 8309 11713 8343 11747
rect 10057 11713 10091 11747
rect 3985 11645 4019 11679
rect 4077 11645 4111 11679
rect 4353 11645 4387 11679
rect 5365 11645 5399 11679
rect 5549 11645 5583 11679
rect 7573 11645 7607 11679
rect 9836 11645 9870 11679
rect 7941 11577 7975 11611
rect 9689 11577 9723 11611
rect 5641 11509 5675 11543
rect 7757 11509 7791 11543
rect 7849 11509 7883 11543
rect 10333 11509 10367 11543
rect 9965 11305 9999 11339
rect 1777 11237 1811 11271
rect 10057 11237 10091 11271
rect 1869 11169 1903 11203
rect 4353 11169 4387 11203
rect 9689 11169 9723 11203
rect 9873 11169 9907 11203
rect 4077 11101 4111 11135
rect 6561 11101 6595 11135
rect 6837 11101 6871 11135
rect 10425 11101 10459 11135
rect 1593 11033 1627 11067
rect 7941 11033 7975 11067
rect 2053 10965 2087 10999
rect 5641 10965 5675 10999
rect 4629 10761 4663 10795
rect 10149 10761 10183 10795
rect 3065 10625 3099 10659
rect 9045 10625 9079 10659
rect 3341 10557 3375 10591
rect 6837 10557 6871 10591
rect 8769 10557 8803 10591
rect 6929 10421 6963 10455
rect 3157 10149 3191 10183
rect 6101 10149 6135 10183
rect 8493 10149 8527 10183
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 4537 10081 4571 10115
rect 4721 10081 4755 10115
rect 5089 10081 5123 10115
rect 6285 10081 6319 10115
rect 7481 10081 7515 10115
rect 4077 10013 4111 10047
rect 4997 10013 5031 10047
rect 2513 9945 2547 9979
rect 7573 9945 7607 9979
rect 8585 10081 8619 10115
rect 10333 10081 10367 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 9873 10013 9907 10047
rect 6377 9877 6411 9911
rect 8493 9877 8527 9911
rect 8677 9877 8711 9911
rect 6285 9673 6319 9707
rect 6561 9673 6595 9707
rect 4721 9537 4755 9571
rect 8769 9537 8803 9571
rect 1869 9469 1903 9503
rect 2053 9469 2087 9503
rect 4997 9469 5031 9503
rect 6469 9469 6503 9503
rect 6561 9469 6595 9503
rect 9321 9469 9355 9503
rect 9597 9469 9631 9503
rect 9781 9469 9815 9503
rect 10701 9469 10735 9503
rect 2421 9401 2455 9435
rect 4905 9401 4939 9435
rect 5457 9401 5491 9435
rect 10793 9333 10827 9367
rect 2973 9129 3007 9163
rect 1685 8993 1719 9027
rect 4261 8993 4295 9027
rect 7849 8993 7883 9027
rect 10333 8993 10367 9027
rect 10517 8993 10551 9027
rect 1409 8925 1443 8959
rect 4445 8789 4479 8823
rect 7941 8789 7975 8823
rect 10609 8789 10643 8823
rect 3617 8585 3651 8619
rect 1593 8517 1627 8551
rect 3617 8449 3651 8483
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 10609 8449 10643 8483
rect 1409 8381 1443 8415
rect 3801 8381 3835 8415
rect 5181 8381 5215 8415
rect 5457 8381 5491 8415
rect 8033 8381 8067 8415
rect 3985 8245 4019 8279
rect 8217 8245 8251 8279
rect 1685 8041 1719 8075
rect 9873 8041 9907 8075
rect 1869 7973 1903 8007
rect 2237 7973 2271 8007
rect 4813 7973 4847 8007
rect 5089 7973 5123 8007
rect 10057 7973 10091 8007
rect 10425 7973 10459 8007
rect 1501 7905 1535 7939
rect 1777 7905 1811 7939
rect 4077 7905 4111 7939
rect 4353 7905 4387 7939
rect 5181 7905 5215 7939
rect 5641 7905 5675 7939
rect 6193 7905 6227 7939
rect 8401 7905 8435 7939
rect 9965 7905 9999 7939
rect 4169 7837 4203 7871
rect 4905 7837 4939 7871
rect 5917 7837 5951 7871
rect 9689 7837 9723 7871
rect 8585 7769 8619 7803
rect 7481 7701 7515 7735
rect 2053 7497 2087 7531
rect 6193 7497 6227 7531
rect 7389 7497 7423 7531
rect 7573 7429 7607 7463
rect 3709 7361 3743 7395
rect 7389 7361 7423 7395
rect 10149 7361 10183 7395
rect 1961 7293 1995 7327
rect 3157 7293 3191 7327
rect 3341 7293 3375 7327
rect 7665 7293 7699 7327
rect 8033 7293 8067 7327
rect 8309 7293 8343 7327
rect 4905 7225 4939 7259
rect 9413 7225 9447 7259
rect 9597 7225 9631 7259
rect 9781 7225 9815 7259
rect 9689 7157 9723 7191
rect 7297 6885 7331 6919
rect 2973 6817 3007 6851
rect 4813 6817 4847 6851
rect 5089 6817 5123 6851
rect 5181 6817 5215 6851
rect 5549 6817 5583 6851
rect 5742 6817 5776 6851
rect 7205 6817 7239 6851
rect 8309 6817 8343 6851
rect 9689 6817 9723 6851
rect 6101 6749 6135 6783
rect 8217 6749 8251 6783
rect 10057 6749 10091 6783
rect 3065 6681 3099 6715
rect 9965 6681 9999 6715
rect 8493 6613 8527 6647
rect 9827 6613 9861 6647
rect 10333 6613 10367 6647
rect 3617 6409 3651 6443
rect 5549 6409 5583 6443
rect 4353 6273 4387 6307
rect 7389 6273 7423 6307
rect 7941 6273 7975 6307
rect 9137 6273 9171 6307
rect 3893 6205 3927 6239
rect 5457 6205 5491 6239
rect 7481 6205 7515 6239
rect 9597 6205 9631 6239
rect 9965 6205 9999 6239
rect 10057 6205 10091 6239
rect 3801 6137 3835 6171
rect 1593 5865 1627 5899
rect 4077 5797 4111 5831
rect 7205 5797 7239 5831
rect 9873 5797 9907 5831
rect 1501 5729 1535 5763
rect 4721 5729 4755 5763
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 6285 5729 6319 5763
rect 6469 5729 6503 5763
rect 6745 5729 6779 5763
rect 8033 5729 8067 5763
rect 8125 5729 8159 5763
rect 8309 5729 8343 5763
rect 9965 5729 9999 5763
rect 4629 5661 4663 5695
rect 8493 5661 8527 5695
rect 6561 5593 6595 5627
rect 6101 5525 6135 5559
rect 9689 5525 9723 5559
rect 10149 5525 10183 5559
rect 1574 5321 1608 5355
rect 3157 5321 3191 5355
rect 5825 5321 5859 5355
rect 1685 5253 1719 5287
rect 7021 5253 7055 5287
rect 9321 5253 9355 5287
rect 1777 5185 1811 5219
rect 4077 5185 4111 5219
rect 4629 5185 4663 5219
rect 1409 5117 1443 5151
rect 2145 5117 2179 5151
rect 3065 5117 3099 5151
rect 4169 5117 4203 5151
rect 5733 5117 5767 5151
rect 6929 5117 6963 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 10609 5117 10643 5151
rect 10793 4981 10827 5015
rect 7297 4777 7331 4811
rect 4077 4709 4111 4743
rect 9873 4709 9907 4743
rect 1593 4641 1627 4675
rect 2145 4641 2179 4675
rect 2329 4641 2363 4675
rect 4261 4641 4295 4675
rect 6009 4641 6043 4675
rect 8217 4641 8251 4675
rect 8401 4641 8435 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 4629 4573 4663 4607
rect 5733 4573 5767 4607
rect 1685 4505 1719 4539
rect 8493 4437 8527 4471
rect 10149 4437 10183 4471
rect 2513 4097 2547 4131
rect 5917 4097 5951 4131
rect 7113 4097 7147 4131
rect 8493 4097 8527 4131
rect 10057 4097 10091 4131
rect 1961 4029 1995 4063
rect 2145 4029 2179 4063
rect 5181 4029 5215 4063
rect 5457 4029 5491 4063
rect 6837 4029 6871 4063
rect 5365 3961 5399 3995
rect 9321 3961 9355 3995
rect 9597 3961 9631 3995
rect 9689 3961 9723 3995
rect 9505 3893 9539 3927
rect 2145 3621 2179 3655
rect 5365 3621 5399 3655
rect 5917 3621 5951 3655
rect 8769 3621 8803 3655
rect 9689 3621 9723 3655
rect 10425 3621 10459 3655
rect 1593 3553 1627 3587
rect 1777 3553 1811 3587
rect 2973 3553 3007 3587
rect 5549 3553 5583 3587
rect 7113 3553 7147 3587
rect 9836 3553 9870 3587
rect 3065 3485 3099 3519
rect 7389 3485 7423 3519
rect 10057 3485 10091 3519
rect 9965 3417 9999 3451
rect 3525 3145 3559 3179
rect 10609 3145 10643 3179
rect 1961 3009 1995 3043
rect 5917 3009 5951 3043
rect 8033 3009 8067 3043
rect 9413 3009 9447 3043
rect 2237 2941 2271 2975
rect 7757 2941 7791 2975
rect 10333 2941 10367 2975
rect 10517 2941 10551 2975
rect 5181 2873 5215 2907
rect 5549 2873 5583 2907
rect 5365 2805 5399 2839
rect 5457 2805 5491 2839
rect 4353 2601 4387 2635
rect 2145 2533 2179 2567
rect 6929 2533 6963 2567
rect 9781 2533 9815 2567
rect 1409 2465 1443 2499
rect 1556 2465 1590 2499
rect 4077 2465 4111 2499
rect 4261 2465 4295 2499
rect 5457 2465 5491 2499
rect 5549 2465 5583 2499
rect 7389 2465 7423 2499
rect 7573 2465 7607 2499
rect 7757 2465 7791 2499
rect 10333 2465 10367 2499
rect 10609 2465 10643 2499
rect 1777 2397 1811 2431
rect 10471 2397 10505 2431
rect 1685 2261 1719 2295
rect 5733 2261 5767 2295
<< metal1 >>
rect 1104 13082 11960 13104
rect 1104 13030 2791 13082
rect 2843 13030 2855 13082
rect 2907 13030 2919 13082
rect 2971 13030 2983 13082
rect 3035 13030 6410 13082
rect 6462 13030 6474 13082
rect 6526 13030 6538 13082
rect 6590 13030 6602 13082
rect 6654 13030 10028 13082
rect 10080 13030 10092 13082
rect 10144 13030 10156 13082
rect 10208 13030 10220 13082
rect 10272 13030 11960 13082
rect 1104 13008 11960 13030
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 9306 12832 9312 12844
rect 4203 12804 9312 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3936 12736 4077 12764
rect 3936 12724 3942 12736
rect 4065 12733 4077 12736
rect 4111 12733 4123 12767
rect 4065 12727 4123 12733
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4304 12736 4353 12764
rect 4304 12724 4310 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4801 12699 4859 12705
rect 4801 12665 4813 12699
rect 4847 12696 4859 12699
rect 5258 12696 5264 12708
rect 4847 12668 5264 12696
rect 4847 12665 4859 12668
rect 4801 12659 4859 12665
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 1104 12538 11960 12560
rect 1104 12486 4600 12538
rect 4652 12486 4664 12538
rect 4716 12486 4728 12538
rect 4780 12486 4792 12538
rect 4844 12486 8219 12538
rect 8271 12486 8283 12538
rect 8335 12486 8347 12538
rect 8399 12486 8411 12538
rect 8463 12486 11960 12538
rect 1104 12464 11960 12486
rect 3878 12316 3884 12368
rect 3936 12356 3942 12368
rect 4338 12356 4344 12368
rect 3936 12328 4344 12356
rect 3936 12316 3942 12328
rect 4338 12316 4344 12328
rect 4396 12316 4402 12368
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2406 12288 2412 12300
rect 2363 12260 2412 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2406 12248 2412 12260
rect 2464 12288 2470 12300
rect 4522 12288 4528 12300
rect 2464 12260 4528 12288
rect 2464 12248 2470 12260
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 5767 12260 5856 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4212 12192 4905 12220
rect 4212 12180 4218 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5408 12192 5457 12220
rect 5408 12180 5414 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5828 12152 5856 12260
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7064 12260 7665 12288
rect 7064 12248 7070 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 8205 12291 8263 12297
rect 8205 12288 8217 12291
rect 7800 12260 8217 12288
rect 7800 12248 7806 12260
rect 8205 12257 8217 12260
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 8665 12223 8723 12229
rect 5960 12192 6005 12220
rect 5960 12180 5966 12192
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 9674 12220 9680 12232
rect 8711 12192 9680 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 5828 12124 7757 12152
rect 7745 12121 7757 12124
rect 7791 12121 7803 12155
rect 7745 12115 7803 12121
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2130 12084 2136 12096
rect 2087 12056 2136 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 6086 12084 6092 12096
rect 2547 12056 6092 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 1104 11994 11960 12016
rect 1104 11942 2791 11994
rect 2843 11942 2855 11994
rect 2907 11942 2919 11994
rect 2971 11942 2983 11994
rect 3035 11942 6410 11994
rect 6462 11942 6474 11994
rect 6526 11942 6538 11994
rect 6590 11942 6602 11994
rect 6654 11942 10028 11994
rect 10080 11942 10092 11994
rect 10144 11942 10156 11994
rect 10208 11942 10220 11994
rect 10272 11942 11960 11994
rect 1104 11920 11960 11942
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 10502 11880 10508 11892
rect 3467 11852 10508 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 5902 11812 5908 11824
rect 3568 11784 4476 11812
rect 3568 11772 3574 11784
rect 4448 11753 4476 11784
rect 5184 11784 5908 11812
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 4982 11744 4988 11756
rect 4479 11716 4988 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 3970 11676 3976 11688
rect 3931 11648 3976 11676
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11676 4399 11679
rect 4522 11676 4528 11688
rect 4387 11648 4528 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 4080 11608 4108 11639
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5184 11608 5212 11784
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 7558 11772 7564 11824
rect 7616 11812 7622 11824
rect 7616 11784 8432 11812
rect 7616 11772 7622 11784
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 5500 11716 8309 11744
rect 5500 11704 5506 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8404 11744 8432 11784
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 9953 11815 10011 11821
rect 9953 11812 9965 11815
rect 9916 11784 9965 11812
rect 9916 11772 9922 11784
rect 9953 11781 9965 11784
rect 9999 11781 10011 11815
rect 9953 11775 10011 11781
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 8404 11716 10057 11744
rect 8297 11707 8355 11713
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 5350 11676 5356 11688
rect 5311 11648 5356 11676
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5534 11676 5540 11688
rect 5495 11648 5540 11676
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 6880 11648 7573 11676
rect 6880 11636 6886 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 9824 11679 9882 11685
rect 9824 11676 9836 11679
rect 7561 11639 7619 11645
rect 7668 11648 9836 11676
rect 4080 11580 5212 11608
rect 5368 11608 5396 11636
rect 7190 11608 7196 11620
rect 5368 11580 7196 11608
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 7668 11608 7696 11648
rect 9824 11645 9836 11648
rect 9870 11645 9882 11679
rect 9824 11639 9882 11645
rect 7926 11608 7932 11620
rect 7300 11580 7696 11608
rect 7887 11580 7932 11608
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 5132 11512 5641 11540
rect 5132 11500 5138 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 7300 11540 7328 11580
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 9674 11608 9680 11620
rect 9587 11580 9680 11608
rect 9674 11568 9680 11580
rect 9732 11608 9738 11620
rect 10686 11608 10692 11620
rect 9732 11580 10692 11608
rect 9732 11568 9738 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 7742 11540 7748 11552
rect 5776 11512 7328 11540
rect 7703 11512 7748 11540
rect 5776 11500 5782 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 8018 11540 8024 11552
rect 7883 11512 8024 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10870 11540 10876 11552
rect 10367 11512 10876 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 1104 11450 11960 11472
rect 1104 11398 4600 11450
rect 4652 11398 4664 11450
rect 4716 11398 4728 11450
rect 4780 11398 4792 11450
rect 4844 11398 8219 11450
rect 8271 11398 8283 11450
rect 8335 11398 8347 11450
rect 8399 11398 8411 11450
rect 8463 11398 11960 11450
rect 1104 11376 11960 11398
rect 3786 11336 3792 11348
rect 1780 11308 3792 11336
rect 1780 11277 1808 11308
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 6178 11336 6184 11348
rect 4028 11308 6184 11336
rect 4028 11296 4034 11308
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 9306 11336 9312 11348
rect 8628 11308 9312 11336
rect 8628 11296 8634 11308
rect 9306 11296 9312 11308
rect 9364 11336 9370 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9364 11308 9965 11336
rect 9364 11296 9370 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11237 1823 11271
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 1765 11231 1823 11237
rect 7484 11240 10057 11268
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 3326 11200 3332 11212
rect 1903 11172 3332 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 3660 11172 4353 11200
rect 3660 11160 3666 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 4982 11160 4988 11212
rect 5040 11200 5046 11212
rect 7484 11200 7512 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 5040 11172 7512 11200
rect 5040 11160 5046 11172
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8076 11172 9689 11200
rect 8076 11160 8082 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3292 11104 4077 11132
rect 3292 11092 3298 11104
rect 4065 11101 4077 11104
rect 4111 11132 4123 11135
rect 6270 11132 6276 11144
rect 4111 11104 6276 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 6270 11092 6276 11104
rect 6328 11132 6334 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6328 11104 6561 11132
rect 6328 11092 6334 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 8110 11132 8116 11144
rect 6871 11104 8116 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9876 11132 9904 11163
rect 10410 11132 10416 11144
rect 9180 11104 9904 11132
rect 10371 11104 10416 11132
rect 9180 11092 9186 11104
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 1627 11036 2728 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 2038 10996 2044 11008
rect 1999 10968 2044 10996
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2700 10996 2728 11036
rect 5460 11036 6592 11064
rect 5460 10996 5488 11036
rect 5626 10996 5632 11008
rect 2700 10968 5488 10996
rect 5587 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6564 10996 6592 11036
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7616 11036 7941 11064
rect 7616 11024 7622 11036
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 6914 10996 6920 11008
rect 6564 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 1104 10906 11960 10928
rect 1104 10854 2791 10906
rect 2843 10854 2855 10906
rect 2907 10854 2919 10906
rect 2971 10854 2983 10906
rect 3035 10854 6410 10906
rect 6462 10854 6474 10906
rect 6526 10854 6538 10906
rect 6590 10854 6602 10906
rect 6654 10854 10028 10906
rect 10080 10854 10092 10906
rect 10144 10854 10156 10906
rect 10208 10854 10220 10906
rect 10272 10854 11960 10906
rect 1104 10832 11960 10854
rect 3786 10752 3792 10804
rect 3844 10792 3850 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 3844 10764 4629 10792
rect 3844 10752 3850 10764
rect 4617 10761 4629 10764
rect 4663 10792 4675 10795
rect 5718 10792 5724 10804
rect 4663 10764 5724 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 9674 10792 9680 10804
rect 7944 10764 9680 10792
rect 7944 10736 7972 10764
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 9732 10764 10149 10792
rect 9732 10752 9738 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 4338 10684 4344 10736
rect 4396 10724 4402 10736
rect 7926 10724 7932 10736
rect 4396 10696 7932 10724
rect 4396 10684 4402 10696
rect 7926 10684 7932 10696
rect 7984 10684 7990 10736
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3234 10656 3240 10668
rect 3099 10628 3240 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 5408 10628 9045 10656
rect 5408 10616 5414 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 4062 10588 4068 10600
rect 3375 10560 4068 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 4948 10560 6837 10588
rect 4948 10548 4954 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 8754 10588 8760 10600
rect 8715 10560 8760 10588
rect 6825 10551 6883 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 6362 10520 6368 10532
rect 6236 10492 6368 10520
rect 6236 10480 6242 10492
rect 6362 10480 6368 10492
rect 6420 10480 6426 10532
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6730 10452 6736 10464
rect 5684 10424 6736 10452
rect 5684 10412 5690 10424
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 9490 10452 9496 10464
rect 6963 10424 9496 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 1104 10362 11960 10384
rect 1104 10310 4600 10362
rect 4652 10310 4664 10362
rect 4716 10310 4728 10362
rect 4780 10310 4792 10362
rect 4844 10310 8219 10362
rect 8271 10310 8283 10362
rect 8335 10310 8347 10362
rect 8399 10310 8411 10362
rect 8463 10310 11960 10362
rect 1104 10288 11960 10310
rect 5534 10248 5540 10260
rect 4540 10220 5540 10248
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 3326 10180 3332 10192
rect 3191 10152 3332 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 1854 10072 1860 10124
rect 1912 10112 1918 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 1912 10084 2421 10112
rect 1912 10072 1918 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3878 10112 3884 10124
rect 2731 10084 3884 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 4540 10121 4568 10220
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 7742 10248 7748 10260
rect 5592 10220 7748 10248
rect 5592 10208 5598 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 5626 10180 5632 10192
rect 4724 10152 5632 10180
rect 4724 10121 4752 10152
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 6086 10180 6092 10192
rect 6047 10152 6092 10180
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 6196 10152 8493 10180
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5994 10112 6000 10124
rect 5123 10084 6000 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 3142 10004 3148 10056
rect 3200 10044 3206 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3200 10016 4077 10044
rect 3200 10004 3206 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4304 10016 4997 10044
rect 4304 10004 4310 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6196 10044 6224 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 10962 10180 10968 10192
rect 8481 10143 8539 10149
rect 10336 10152 10968 10180
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10112 6331 10115
rect 6362 10112 6368 10124
rect 6319 10084 6368 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 7466 10112 7472 10124
rect 7427 10084 7472 10112
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9306 10112 9312 10124
rect 8619 10084 9312 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10336 10121 10364 10152
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 10870 10112 10876 10124
rect 10735 10084 10876 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 6144 10016 6224 10044
rect 6380 10044 6408 10072
rect 9214 10044 9220 10056
rect 6380 10016 9220 10044
rect 6144 10004 6150 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9824 10016 9873 10044
rect 9824 10004 9830 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 2498 9976 2504 9988
rect 2459 9948 2504 9976
rect 2498 9936 2504 9948
rect 2556 9936 2562 9988
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 5000 9948 7573 9976
rect 5000 9920 5028 9948
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 10520 9976 10548 10075
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 7561 9939 7619 9945
rect 7668 9948 10548 9976
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4706 9908 4712 9920
rect 4396 9880 4712 9908
rect 4396 9868 4402 9880
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 4982 9868 4988 9920
rect 5040 9868 5046 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 5592 9880 6377 9908
rect 5592 9868 5598 9880
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 7668 9908 7696 9948
rect 6788 9880 7696 9908
rect 8481 9911 8539 9917
rect 6788 9868 6794 9880
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 8527 9880 8677 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 8665 9877 8677 9880
rect 8711 9908 8723 9911
rect 8938 9908 8944 9920
rect 8711 9880 8944 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 1104 9818 11960 9840
rect 1104 9766 2791 9818
rect 2843 9766 2855 9818
rect 2907 9766 2919 9818
rect 2971 9766 2983 9818
rect 3035 9766 6410 9818
rect 6462 9766 6474 9818
rect 6526 9766 6538 9818
rect 6590 9766 6602 9818
rect 6654 9766 10028 9818
rect 10080 9766 10092 9818
rect 10144 9766 10156 9818
rect 10208 9766 10220 9818
rect 10272 9766 11960 9818
rect 1104 9744 11960 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 6086 9704 6092 9716
rect 1912 9676 6092 9704
rect 1912 9664 1918 9676
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 6270 9704 6276 9716
rect 6183 9676 6276 9704
rect 6270 9664 6276 9676
rect 6328 9704 6334 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 6328 9676 6561 9704
rect 6328 9664 6334 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 10410 9636 10416 9648
rect 1872 9608 10416 9636
rect 1872 9509 1900 9608
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5166 9568 5172 9580
rect 4755 9540 5172 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 6052 9540 8769 9568
rect 6052 9528 6058 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9214 9528 9220 9580
rect 9272 9568 9278 9580
rect 9272 9540 10732 9568
rect 9272 9528 9278 9540
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 4985 9503 5043 9509
rect 2087 9472 4292 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9401 2467 9435
rect 2409 9395 2467 9401
rect 2424 9364 2452 9395
rect 3970 9364 3976 9376
rect 2424 9336 3976 9364
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4264 9364 4292 9472
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5534 9500 5540 9512
rect 5031 9472 5540 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6086 9500 6092 9512
rect 5868 9472 6092 9500
rect 5868 9460 5874 9472
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 6236 9472 6469 9500
rect 6236 9460 6242 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9500 6607 9503
rect 8662 9500 8668 9512
rect 6595 9472 8668 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 9180 9472 9321 9500
rect 9180 9460 9186 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4396 9404 4905 9432
rect 4396 9392 4402 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 4893 9395 4951 9401
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 6730 9432 6736 9444
rect 5491 9404 6736 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 9600 9432 9628 9463
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10704 9509 10732 9540
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9732 9472 9781 9500
rect 9732 9460 9738 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 7984 9404 9628 9432
rect 7984 9392 7990 9404
rect 10318 9364 10324 9376
rect 4264 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 10468 9336 10793 9364
rect 10468 9324 10474 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 1104 9274 11960 9296
rect 1104 9222 4600 9274
rect 4652 9222 4664 9274
rect 4716 9222 4728 9274
rect 4780 9222 4792 9274
rect 4844 9222 8219 9274
rect 8271 9222 8283 9274
rect 8335 9222 8347 9274
rect 8399 9222 8411 9274
rect 8463 9222 11960 9274
rect 1104 9200 11960 9222
rect 2958 9160 2964 9172
rect 2871 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9160 3022 9172
rect 4246 9160 4252 9172
rect 3016 9132 4252 9160
rect 3016 9120 3022 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 3936 9064 7420 9092
rect 3936 9052 3942 9064
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 3896 9024 3924 9052
rect 7392 9036 7420 9064
rect 2372 8996 3924 9024
rect 4249 9027 4307 9033
rect 2372 8984 2378 8996
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 5534 9024 5540 9036
rect 4295 8996 5540 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7432 8996 7849 9024
rect 7432 8984 7438 8996
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 7837 8987 7895 8993
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 10410 9024 10416 9036
rect 10367 8996 10416 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 3234 8956 3240 8968
rect 1397 8919 1455 8925
rect 2332 8928 3240 8956
rect 1412 8820 1440 8919
rect 2332 8820 2360 8928
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 5994 8956 6000 8968
rect 4028 8928 6000 8956
rect 4028 8916 4034 8928
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 10520 8956 10548 8987
rect 9456 8928 10548 8956
rect 9456 8916 9462 8928
rect 2958 8848 2964 8900
rect 3016 8848 3022 8900
rect 1412 8792 2360 8820
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 2976 8820 3004 8848
rect 2740 8792 3004 8820
rect 2740 8780 2746 8792
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 4304 8792 4445 8820
rect 4304 8780 4310 8792
rect 4433 8789 4445 8792
rect 4479 8789 4491 8823
rect 4433 8783 4491 8789
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 7006 8820 7012 8832
rect 4580 8792 7012 8820
rect 4580 8780 4586 8792
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7340 8792 7941 8820
rect 7340 8780 7346 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 10594 8820 10600 8832
rect 10555 8792 10600 8820
rect 7929 8783 7987 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 1104 8730 11960 8752
rect 1104 8678 2791 8730
rect 2843 8678 2855 8730
rect 2907 8678 2919 8730
rect 2971 8678 2983 8730
rect 3035 8678 6410 8730
rect 6462 8678 6474 8730
rect 6526 8678 6538 8730
rect 6590 8678 6602 8730
rect 6654 8678 10028 8730
rect 10080 8678 10092 8730
rect 10144 8678 10156 8730
rect 10208 8678 10220 8730
rect 10272 8678 11960 8730
rect 1104 8656 11960 8678
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 9122 8616 9128 8628
rect 3651 8588 9128 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8548 1642 8560
rect 6822 8548 6828 8560
rect 1636 8520 6828 8548
rect 1636 8508 1642 8520
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4522 8480 4528 8492
rect 3651 8452 3832 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8412 1458 8424
rect 3694 8412 3700 8424
rect 1452 8384 3700 8412
rect 1452 8372 1458 8384
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 3804 8421 3832 8452
rect 3896 8452 4528 8480
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3896 8344 3924 8452
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5718 8480 5724 8492
rect 5307 8452 5724 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7466 8480 7472 8492
rect 5951 8452 7472 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8812 8452 9229 8480
rect 8812 8440 8818 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9490 8480 9496 8492
rect 9451 8452 9496 8480
rect 9217 8443 9275 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 9640 8452 10609 8480
rect 9640 8440 9646 8452
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4028 8384 5181 8412
rect 4028 8372 4034 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 5169 8375 5227 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5736 8412 5764 8440
rect 6086 8412 6092 8424
rect 5736 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 9858 8412 9864 8424
rect 9180 8384 9864 8412
rect 9180 8372 9186 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 3896 8316 4016 8344
rect 3988 8285 4016 8316
rect 5460 8316 8248 8344
rect 5460 8288 5488 8316
rect 3973 8279 4031 8285
rect 3973 8245 3985 8279
rect 4019 8245 4031 8279
rect 3973 8239 4031 8245
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5442 8276 5448 8288
rect 5224 8248 5448 8276
rect 5224 8236 5230 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 8220 8285 8248 8316
rect 8205 8279 8263 8285
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8570 8276 8576 8288
rect 8251 8248 8576 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 1104 8186 11960 8208
rect 1104 8134 4600 8186
rect 4652 8134 4664 8186
rect 4716 8134 4728 8186
rect 4780 8134 4792 8186
rect 4844 8134 8219 8186
rect 8271 8134 8283 8186
rect 8335 8134 8347 8186
rect 8399 8134 8411 8186
rect 8463 8134 11960 8186
rect 1104 8112 11960 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 2498 8072 2504 8084
rect 1719 8044 2504 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 7650 8072 7656 8084
rect 4632 8044 7656 8072
rect 4632 8016 4660 8044
rect 7650 8032 7656 8044
rect 7708 8072 7714 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 7708 8044 9873 8072
rect 7708 8032 7714 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 1854 8004 1860 8016
rect 1815 7976 1860 8004
rect 1854 7964 1860 7976
rect 1912 7964 1918 8016
rect 2225 8007 2283 8013
rect 2225 7973 2237 8007
rect 2271 8004 2283 8007
rect 3602 8004 3608 8016
rect 2271 7976 3608 8004
rect 2271 7973 2283 7976
rect 2225 7967 2283 7973
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4614 7964 4620 8016
rect 4672 7964 4678 8016
rect 4801 8007 4859 8013
rect 4801 7973 4813 8007
rect 4847 8004 4859 8007
rect 4890 8004 4896 8016
rect 4847 7976 4896 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 5074 8004 5080 8016
rect 5035 7976 5080 8004
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 8202 8004 8208 8016
rect 7064 7976 8208 8004
rect 7064 7964 7070 7976
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 10045 8007 10103 8013
rect 10045 8004 10057 8007
rect 8812 7976 10057 8004
rect 8812 7964 8818 7976
rect 10045 7973 10057 7976
rect 10091 7973 10103 8007
rect 10045 7967 10103 7973
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 10413 8007 10471 8013
rect 10413 8004 10425 8007
rect 10376 7976 10425 8004
rect 10376 7964 10382 7976
rect 10413 7973 10425 7976
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 1489 7939 1547 7945
rect 1489 7936 1501 7939
rect 1412 7908 1501 7936
rect 1412 7732 1440 7908
rect 1489 7905 1501 7908
rect 1535 7905 1547 7939
rect 1489 7899 1547 7905
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2038 7936 2044 7948
rect 1811 7908 2044 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2038 7896 2044 7908
rect 2096 7936 2102 7948
rect 4065 7939 4123 7945
rect 2096 7908 4016 7936
rect 2096 7896 2102 7908
rect 3988 7800 4016 7908
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4246 7936 4252 7948
rect 4111 7908 4252 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4246 7896 4252 7908
rect 4304 7896 4310 7948
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 4522 7936 4528 7948
rect 4387 7908 4528 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 5675 7908 6193 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 6972 7908 8401 7936
rect 6972 7896 6978 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 4154 7868 4160 7880
rect 4115 7840 4160 7868
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4890 7868 4896 7880
rect 4803 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7868 4954 7880
rect 5442 7868 5448 7880
rect 4948 7840 5448 7868
rect 4948 7828 4954 7840
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6270 7868 6276 7880
rect 5951 7840 6276 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 6880 7840 9689 7868
rect 6880 7828 6886 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9968 7868 9996 7899
rect 9677 7831 9735 7837
rect 9876 7840 9996 7868
rect 5074 7800 5080 7812
rect 3988 7772 5080 7800
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 8018 7800 8024 7812
rect 7708 7772 8024 7800
rect 7708 7760 7714 7772
rect 8018 7760 8024 7772
rect 8076 7800 8082 7812
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 8076 7772 8585 7800
rect 8076 7760 8082 7772
rect 8573 7769 8585 7772
rect 8619 7800 8631 7803
rect 9876 7800 9904 7840
rect 8619 7772 9904 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 4154 7732 4160 7744
rect 1412 7704 4160 7732
rect 4154 7692 4160 7704
rect 4212 7732 4218 7744
rect 7282 7732 7288 7744
rect 4212 7704 7288 7732
rect 4212 7692 4218 7704
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 7742 7732 7748 7744
rect 7515 7704 7748 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 1104 7642 11960 7664
rect 1104 7590 2791 7642
rect 2843 7590 2855 7642
rect 2907 7590 2919 7642
rect 2971 7590 2983 7642
rect 3035 7590 6410 7642
rect 6462 7590 6474 7642
rect 6526 7590 6538 7642
rect 6590 7590 6602 7642
rect 6654 7590 10028 7642
rect 10080 7590 10092 7642
rect 10144 7590 10156 7642
rect 10208 7590 10220 7642
rect 10272 7590 11960 7642
rect 1104 7568 11960 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2130 7528 2136 7540
rect 2087 7500 2136 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2130 7488 2136 7500
rect 2188 7528 2194 7540
rect 2590 7528 2596 7540
rect 2188 7500 2596 7528
rect 2188 7488 2194 7500
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 6178 7528 6184 7540
rect 6139 7500 6184 7528
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7528 7435 7531
rect 9490 7528 9496 7540
rect 7423 7500 9496 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 4304 7432 7573 7460
rect 4304 7420 4310 7432
rect 7561 7429 7573 7432
rect 7607 7429 7619 7463
rect 7561 7423 7619 7429
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 8168 7432 10180 7460
rect 8168 7420 8174 7432
rect 3697 7395 3755 7401
rect 1964 7364 3648 7392
rect 1964 7333 1992 7364
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7293 2007 7327
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 1949 7287 2007 7293
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3418 7324 3424 7336
rect 3375 7296 3424 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3620 7324 3648 7364
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 5166 7392 5172 7404
rect 3743 7364 5172 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 5500 7364 7389 7392
rect 5500 7352 5506 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 9582 7392 9588 7404
rect 7377 7355 7435 7361
rect 7668 7364 9588 7392
rect 5718 7324 5724 7336
rect 3620 7296 5724 7324
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 7466 7324 7472 7336
rect 7340 7296 7472 7324
rect 7340 7284 7346 7296
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 7668 7333 7696 7364
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 10152 7401 10180 7432
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 8018 7324 8024 7336
rect 7979 7296 8024 7324
rect 7653 7287 7711 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 3292 7228 4905 7256
rect 3292 7216 3298 7228
rect 4893 7225 4905 7228
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 8312 7256 8340 7287
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9364 7296 9812 7324
rect 9364 7284 9370 7296
rect 7248 7228 8340 7256
rect 9401 7259 9459 7265
rect 7248 7216 7254 7228
rect 9401 7225 9413 7259
rect 9447 7225 9459 7259
rect 9401 7219 9459 7225
rect 2498 7148 2504 7200
rect 2556 7188 2562 7200
rect 3510 7188 3516 7200
rect 2556 7160 3516 7188
rect 2556 7148 2562 7160
rect 3510 7148 3516 7160
rect 3568 7188 3574 7200
rect 5442 7188 5448 7200
rect 3568 7160 5448 7188
rect 3568 7148 3574 7160
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 7374 7188 7380 7200
rect 6328 7160 7380 7188
rect 6328 7148 6334 7160
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 9416 7188 9444 7219
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 9784 7265 9812 7296
rect 9585 7259 9643 7265
rect 9585 7256 9597 7259
rect 9548 7228 9597 7256
rect 9548 7216 9554 7228
rect 9585 7225 9597 7228
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 9674 7188 9680 7200
rect 7524 7160 9444 7188
rect 9635 7160 9680 7188
rect 7524 7148 7530 7160
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 1104 7098 11960 7120
rect 1104 7046 4600 7098
rect 4652 7046 4664 7098
rect 4716 7046 4728 7098
rect 4780 7046 4792 7098
rect 4844 7046 8219 7098
rect 8271 7046 8283 7098
rect 8335 7046 8347 7098
rect 8399 7046 8411 7098
rect 8463 7046 11960 7098
rect 1104 7024 11960 7046
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 9674 6984 9680 6996
rect 5132 6956 9680 6984
rect 5132 6944 5138 6956
rect 9674 6944 9680 6956
rect 9732 6984 9738 6996
rect 10778 6984 10784 6996
rect 9732 6956 10784 6984
rect 9732 6944 9738 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 5442 6916 5448 6928
rect 5092 6888 5448 6916
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 2976 6780 3004 6811
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 3602 6848 3608 6860
rect 3200 6820 3608 6848
rect 3200 6808 3206 6820
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 5092 6857 5120 6888
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 6270 6916 6276 6928
rect 5552 6888 6276 6916
rect 5552 6857 5580 6888
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 7282 6916 7288 6928
rect 7243 6888 7288 6916
rect 7282 6876 7288 6888
rect 7340 6876 7346 6928
rect 9600 6888 9812 6916
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4212 6820 4813 6848
rect 4212 6808 4218 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 2976 6752 3924 6780
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3786 6712 3792 6724
rect 3099 6684 3792 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3786 6672 3792 6684
rect 3844 6672 3850 6724
rect 3896 6712 3924 6752
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 5184 6780 5212 6811
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5730 6851 5788 6857
rect 5730 6848 5742 6851
rect 5684 6820 5742 6848
rect 5684 6808 5690 6820
rect 5730 6817 5742 6820
rect 5776 6817 5788 6851
rect 5730 6811 5788 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 7156 6820 7205 6848
rect 7156 6808 7162 6820
rect 7193 6817 7205 6820
rect 7239 6817 7251 6851
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 7193 6811 7251 6817
rect 7392 6820 8309 6848
rect 4304 6752 5212 6780
rect 4304 6740 4310 6752
rect 4614 6712 4620 6724
rect 3896 6684 4620 6712
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 5184 6712 5212 6752
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5316 6752 6101 6780
rect 5316 6740 5322 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7392 6780 7420 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 6880 6752 7420 6780
rect 7484 6752 8217 6780
rect 6880 6740 6886 6752
rect 5442 6712 5448 6724
rect 5184 6684 5448 6712
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 6270 6672 6276 6724
rect 6328 6712 6334 6724
rect 7484 6712 7512 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 9600 6780 9628 6888
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9784 6848 9812 6888
rect 9784 6820 10088 6848
rect 9677 6811 9735 6817
rect 8205 6743 8263 6749
rect 8312 6752 9628 6780
rect 6328 6684 7512 6712
rect 6328 6672 6334 6684
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8312 6712 8340 6752
rect 9692 6712 9720 6811
rect 10060 6789 10088 6820
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 9950 6712 9956 6724
rect 8168 6684 8340 6712
rect 8404 6684 9720 6712
rect 9911 6684 9956 6712
rect 8168 6672 8174 6684
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 8404 6644 8432 6684
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 3476 6616 8432 6644
rect 3476 6604 3482 6616
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8536 6616 8581 6644
rect 8536 6604 8542 6616
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9815 6647 9873 6653
rect 9815 6644 9827 6647
rect 9732 6616 9827 6644
rect 9732 6604 9738 6616
rect 9815 6613 9827 6616
rect 9861 6613 9873 6647
rect 10318 6644 10324 6656
rect 10279 6616 10324 6644
rect 9815 6607 9873 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 1104 6554 11960 6576
rect 1104 6502 2791 6554
rect 2843 6502 2855 6554
rect 2907 6502 2919 6554
rect 2971 6502 2983 6554
rect 3035 6502 6410 6554
rect 6462 6502 6474 6554
rect 6526 6502 6538 6554
rect 6590 6502 6602 6554
rect 6654 6502 10028 6554
rect 10080 6502 10092 6554
rect 10144 6502 10156 6554
rect 10208 6502 10220 6554
rect 10272 6502 11960 6554
rect 1104 6480 11960 6502
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 4890 6440 4896 6452
rect 3651 6412 4896 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 8478 6440 8484 6452
rect 5776 6412 8484 6440
rect 5776 6400 5782 6412
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 3878 6372 3884 6384
rect 3620 6344 3884 6372
rect 3620 6168 3648 6344
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 5350 6372 5356 6384
rect 4356 6344 5356 6372
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4356 6313 4384 6344
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 5442 6332 5448 6384
rect 5500 6372 5506 6384
rect 9306 6372 9312 6384
rect 5500 6344 9312 6372
rect 5500 6332 5506 6344
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 10502 6372 10508 6384
rect 10008 6344 10508 6372
rect 10008 6332 10014 6344
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 4341 6307 4399 6313
rect 3752 6276 4292 6304
rect 3752 6264 3758 6276
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 3789 6171 3847 6177
rect 3789 6168 3801 6171
rect 3620 6140 3801 6168
rect 3789 6137 3801 6140
rect 3835 6137 3847 6171
rect 4264 6168 4292 6276
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6822 6304 6828 6316
rect 5592 6276 6828 6304
rect 5592 6264 5598 6276
rect 6822 6264 6828 6276
rect 6880 6304 6886 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6880 6276 7389 6304
rect 6880 6264 6886 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7926 6304 7932 6316
rect 7616 6276 7696 6304
rect 7887 6276 7932 6304
rect 7616 6264 7622 6276
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5350 6236 5356 6248
rect 4856 6208 5356 6236
rect 4856 6196 4862 6208
rect 5350 6196 5356 6208
rect 5408 6236 5414 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5408 6208 5457 6236
rect 5408 6196 5414 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7524 6208 7569 6236
rect 7524 6196 7530 6208
rect 5810 6168 5816 6180
rect 4264 6140 5816 6168
rect 3789 6131 3847 6137
rect 5810 6128 5816 6140
rect 5868 6168 5874 6180
rect 6270 6168 6276 6180
rect 5868 6140 6276 6168
rect 5868 6128 5874 6140
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 7668 6168 7696 6276
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9214 6304 9220 6316
rect 9171 6276 9220 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8018 6236 8024 6248
rect 7800 6208 8024 6236
rect 7800 6196 7806 6208
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6236 10103 6239
rect 10502 6236 10508 6248
rect 10091 6208 10508 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 7926 6168 7932 6180
rect 7668 6140 7932 6168
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3602 6100 3608 6112
rect 2740 6072 3608 6100
rect 2740 6060 2746 6072
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 7558 6100 7564 6112
rect 3752 6072 7564 6100
rect 3752 6060 3758 6072
rect 7558 6060 7564 6072
rect 7616 6100 7622 6112
rect 9968 6100 9996 6199
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 7616 6072 9996 6100
rect 7616 6060 7622 6072
rect 1104 6010 11960 6032
rect 1104 5958 4600 6010
rect 4652 5958 4664 6010
rect 4716 5958 4728 6010
rect 4780 5958 4792 6010
rect 4844 5958 8219 6010
rect 8271 5958 8283 6010
rect 8335 5958 8347 6010
rect 8399 5958 8411 6010
rect 8463 5958 11960 6010
rect 1104 5936 11960 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 3142 5896 3148 5908
rect 1627 5868 3148 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3660 5868 8340 5896
rect 3660 5856 3666 5868
rect 4062 5828 4068 5840
rect 4023 5800 4068 5828
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 7193 5831 7251 5837
rect 4212 5800 6868 5828
rect 4212 5788 4218 5800
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 2222 5760 2228 5772
rect 1535 5732 2228 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 4246 5760 4252 5772
rect 3752 5732 4252 5760
rect 3752 5720 3758 5732
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5760 4767 5763
rect 4982 5760 4988 5772
rect 4755 5732 4988 5760
rect 4755 5729 4767 5732
rect 4709 5723 4767 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 5258 5760 5264 5772
rect 5132 5732 5177 5760
rect 5219 5732 5264 5760
rect 5132 5720 5138 5732
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6472 5769 6500 5800
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6236 5732 6285 5760
rect 6236 5720 6242 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6273 5723 6331 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6604 5732 6745 5760
rect 6604 5720 6610 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6840 5760 6868 5800
rect 7193 5797 7205 5831
rect 7239 5828 7251 5831
rect 7466 5828 7472 5840
rect 7239 5800 7472 5828
rect 7239 5797 7251 5800
rect 7193 5791 7251 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 8202 5828 8208 5840
rect 7576 5800 8208 5828
rect 7576 5760 7604 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 6840 5732 7604 5760
rect 6733 5723 6791 5729
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7984 5732 8033 5760
rect 7984 5720 7990 5732
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8312 5769 8340 5868
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8754 5828 8760 5840
rect 8444 5800 8760 5828
rect 8444 5788 8450 5800
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 9861 5831 9919 5837
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 10594 5828 10600 5840
rect 9907 5800 10600 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 8297 5763 8355 5769
rect 8168 5732 8213 5760
rect 8168 5720 8174 5732
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 9306 5760 9312 5772
rect 8343 5732 9312 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9950 5760 9956 5772
rect 9911 5732 9956 5760
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 3200 5664 4629 5692
rect 3200 5652 3206 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 4617 5655 4675 5661
rect 5644 5664 8493 5692
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 2406 5624 2412 5636
rect 1452 5596 2412 5624
rect 1452 5584 1458 5596
rect 2406 5584 2412 5596
rect 2464 5624 2470 5636
rect 5644 5624 5672 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9214 5692 9220 5704
rect 8720 5664 9220 5692
rect 8720 5652 8726 5664
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 2464 5596 5672 5624
rect 6549 5627 6607 5633
rect 2464 5584 2470 5596
rect 6549 5593 6561 5627
rect 6595 5624 6607 5627
rect 7282 5624 7288 5636
rect 6595 5596 7288 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 7282 5584 7288 5596
rect 7340 5624 7346 5636
rect 8110 5624 8116 5636
rect 7340 5596 8116 5624
rect 7340 5584 7346 5596
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 8220 5596 10180 5624
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6822 5556 6828 5568
rect 6135 5528 6828 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8220 5556 8248 5596
rect 8076 5528 8248 5556
rect 8076 5516 8082 5528
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9490 5556 9496 5568
rect 8628 5528 9496 5556
rect 8628 5516 8634 5528
rect 9490 5516 9496 5528
rect 9548 5556 9554 5568
rect 10152 5565 10180 5596
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9548 5528 9689 5556
rect 9548 5516 9554 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 9677 5519 9735 5525
rect 10137 5559 10195 5565
rect 10137 5525 10149 5559
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 1104 5466 11960 5488
rect 1104 5414 2791 5466
rect 2843 5414 2855 5466
rect 2907 5414 2919 5466
rect 2971 5414 2983 5466
rect 3035 5414 6410 5466
rect 6462 5414 6474 5466
rect 6526 5414 6538 5466
rect 6590 5414 6602 5466
rect 6654 5414 10028 5466
rect 10080 5414 10092 5466
rect 10144 5414 10156 5466
rect 10208 5414 10220 5466
rect 10272 5414 11960 5466
rect 1104 5392 11960 5414
rect 1562 5355 1620 5361
rect 1562 5321 1574 5355
rect 1608 5352 1620 5355
rect 3145 5355 3203 5361
rect 1608 5324 3096 5352
rect 1608 5321 1620 5324
rect 1562 5315 1620 5321
rect 1670 5284 1676 5296
rect 1631 5256 1676 5284
rect 1670 5244 1676 5256
rect 1728 5244 1734 5296
rect 3068 5284 3096 5324
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3878 5352 3884 5364
rect 3191 5324 3884 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 7190 5352 7196 5364
rect 5859 5324 7196 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 7190 5312 7196 5324
rect 7248 5352 7254 5364
rect 9582 5352 9588 5364
rect 7248 5324 9588 5352
rect 7248 5312 7254 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 5718 5284 5724 5296
rect 3068 5256 5724 5284
rect 5718 5244 5724 5256
rect 5776 5284 5782 5296
rect 6270 5284 6276 5296
rect 5776 5256 6276 5284
rect 5776 5244 5782 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 6972 5256 7021 5284
rect 6972 5244 6978 5256
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9309 5287 9367 5293
rect 9309 5284 9321 5287
rect 9180 5256 9321 5284
rect 9180 5244 9186 5256
rect 9309 5253 9321 5256
rect 9355 5253 9367 5287
rect 9309 5247 9367 5253
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3844 5188 4077 5216
rect 3844 5176 3850 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 9674 5216 9680 5228
rect 4663 5188 9680 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 2130 5148 2136 5160
rect 2091 5120 2136 5148
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3326 5148 3332 5160
rect 3099 5120 3332 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 5166 5148 5172 5160
rect 4203 5120 5172 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6638 5148 6644 5160
rect 5767 5120 6644 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8662 5148 8668 5160
rect 8251 5120 8668 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7944 5080 7972 5111
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 10594 5148 10600 5160
rect 10555 5120 10600 5148
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 6880 5052 7972 5080
rect 6880 5040 6886 5052
rect 9582 5040 9588 5092
rect 9640 5080 9646 5092
rect 10870 5080 10876 5092
rect 9640 5052 10876 5080
rect 9640 5040 9646 5052
rect 10870 5040 10876 5052
rect 10928 5040 10934 5092
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 9272 4984 10793 5012
rect 9272 4972 9278 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 1104 4922 11960 4944
rect 1104 4870 4600 4922
rect 4652 4870 4664 4922
rect 4716 4870 4728 4922
rect 4780 4870 4792 4922
rect 4844 4870 8219 4922
rect 8271 4870 8283 4922
rect 8335 4870 8347 4922
rect 8399 4870 8411 4922
rect 8463 4870 11960 4922
rect 1104 4848 11960 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1820 4780 5672 4808
rect 1820 4768 1826 4780
rect 1670 4740 1676 4752
rect 1583 4712 1676 4740
rect 1596 4681 1624 4712
rect 1670 4700 1676 4712
rect 1728 4740 1734 4752
rect 4065 4743 4123 4749
rect 1728 4712 2544 4740
rect 1728 4700 1734 4712
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4641 2191 4675
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2133 4635 2191 4641
rect 2148 4604 2176 4635
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2516 4604 2544 4712
rect 4065 4709 4077 4743
rect 4111 4740 4123 4743
rect 4154 4740 4160 4752
rect 4111 4712 4160 4740
rect 4111 4709 4123 4712
rect 4065 4703 4123 4709
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 5644 4740 5672 4780
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 7282 4808 7288 4820
rect 6328 4780 6684 4808
rect 7243 4780 7288 4808
rect 6328 4768 6334 4780
rect 6656 4740 6684 4780
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 10594 4808 10600 4820
rect 9692 4780 10600 4808
rect 9692 4740 9720 4780
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 5644 4712 5856 4740
rect 6656 4712 9720 4740
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 3786 4672 3792 4684
rect 3660 4644 3792 4672
rect 3660 4632 3666 4644
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4890 4672 4896 4684
rect 4295 4644 4896 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 2148 4576 2268 4604
rect 2516 4576 4629 4604
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4505 1731 4539
rect 2240 4536 2268 4576
rect 4617 4573 4629 4576
rect 4663 4604 4675 4607
rect 5534 4604 5540 4616
rect 4663 4576 5540 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5828 4604 5856 4712
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9824 4712 9873 4740
rect 9824 4700 9830 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 7742 4672 7748 4684
rect 6104 4644 7748 4672
rect 6104 4604 6132 4644
rect 7742 4632 7748 4644
rect 7800 4672 7806 4684
rect 8202 4672 8208 4684
rect 7800 4644 8208 4672
rect 7800 4632 7806 4644
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 5828 4576 6132 4604
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 7926 4604 7932 4616
rect 6236 4576 7932 4604
rect 6236 4564 6242 4576
rect 7926 4564 7932 4576
rect 7984 4604 7990 4616
rect 8404 4604 8432 4635
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9548 4644 9689 4672
rect 9548 4632 9554 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10318 4672 10324 4684
rect 9999 4644 10324 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 7984 4576 8432 4604
rect 7984 4564 7990 4576
rect 4982 4536 4988 4548
rect 2240 4508 4988 4536
rect 1673 4499 1731 4505
rect 1688 4468 1716 4499
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 9030 4536 9036 4548
rect 7668 4508 9036 4536
rect 3970 4468 3976 4480
rect 1688 4440 3976 4468
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 7668 4468 7696 4508
rect 9030 4496 9036 4508
rect 9088 4496 9094 4548
rect 5316 4440 7696 4468
rect 5316 4428 5322 4440
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 7800 4440 8493 4468
rect 7800 4428 7806 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 9582 4468 9588 4480
rect 8720 4440 9588 4468
rect 8720 4428 8726 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 9824 4440 10149 4468
rect 9824 4428 9830 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 1104 4378 11960 4400
rect 1104 4326 2791 4378
rect 2843 4326 2855 4378
rect 2907 4326 2919 4378
rect 2971 4326 2983 4378
rect 3035 4326 6410 4378
rect 6462 4326 6474 4378
rect 6526 4326 6538 4378
rect 6590 4326 6602 4378
rect 6654 4326 10028 4378
rect 10080 4326 10092 4378
rect 10144 4326 10156 4378
rect 10208 4326 10220 4378
rect 10272 4326 11960 4378
rect 1104 4304 11960 4326
rect 2148 4236 4108 4264
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2148 4069 2176 4236
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 4080 4196 4108 4236
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 9490 4264 9496 4276
rect 7064 4236 9496 4264
rect 7064 4224 7070 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 6178 4196 6184 4208
rect 2648 4168 3556 4196
rect 4080 4168 6184 4196
rect 2648 4156 2654 4168
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 3418 4128 3424 4140
rect 2547 4100 3424 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3528 4128 3556 4168
rect 6178 4156 6184 4168
rect 6236 4156 6242 4208
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 8202 4196 8208 4208
rect 7984 4168 8208 4196
rect 7984 4156 7990 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 9214 4196 9220 4208
rect 8312 4168 9220 4196
rect 5902 4128 5908 4140
rect 3528 4100 5212 4128
rect 5863 4100 5908 4128
rect 5184 4072 5212 4100
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 6788 4100 7113 4128
rect 6788 4088 6794 4100
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 8312 4128 8340 4168
rect 9214 4156 9220 4168
rect 9272 4156 9278 4208
rect 7248 4100 8340 4128
rect 8481 4131 8539 4137
rect 7248 4088 7254 4100
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8846 4128 8852 4140
rect 8527 4100 8852 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9640 4100 10057 4128
rect 9640 4088 9646 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 5166 4060 5172 4072
rect 2372 4032 4108 4060
rect 5127 4032 5172 4060
rect 2372 4020 2378 4032
rect 4080 3992 4108 4032
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5442 4060 5448 4072
rect 5403 4032 5448 4060
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6822 4060 6828 4072
rect 5776 4032 6828 4060
rect 5776 4020 5782 4032
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7432 4032 7788 4060
rect 7432 4020 7438 4032
rect 5353 3995 5411 4001
rect 5353 3992 5365 3995
rect 4080 3964 5365 3992
rect 5353 3961 5365 3964
rect 5399 3961 5411 3995
rect 7760 3992 7788 4032
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 8996 4032 9628 4060
rect 8996 4020 9002 4032
rect 9600 4001 9628 4032
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 7760 3964 9321 3992
rect 5353 3955 5411 3961
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3961 9643 3995
rect 9585 3955 9643 3961
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 10778 3992 10784 4004
rect 9723 3964 10784 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 5684 3896 9505 3924
rect 5684 3884 5690 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 1104 3834 11960 3856
rect 1104 3782 4600 3834
rect 4652 3782 4664 3834
rect 4716 3782 4728 3834
rect 4780 3782 4792 3834
rect 4844 3782 8219 3834
rect 8271 3782 8283 3834
rect 8335 3782 8347 3834
rect 8399 3782 8411 3834
rect 8463 3782 11960 3834
rect 1104 3760 11960 3782
rect 4246 3720 4252 3732
rect 1559 3692 4252 3720
rect 1559 3593 1587 3692
rect 4246 3680 4252 3692
rect 4304 3720 4310 3732
rect 5074 3720 5080 3732
rect 4304 3692 5080 3720
rect 4304 3680 4310 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5592 3692 9720 3720
rect 5592 3680 5598 3692
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2314 3652 2320 3664
rect 2179 3624 2320 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 5350 3652 5356 3664
rect 5311 3624 5356 3652
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 5718 3652 5724 3664
rect 5460 3624 5724 3652
rect 1559 3587 1639 3593
rect 1559 3556 1593 3587
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1581 3547 1639 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3510 3584 3516 3596
rect 3007 3556 3516 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 5460 3584 5488 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 6086 3652 6092 3664
rect 5951 3624 6092 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 8754 3652 8760 3664
rect 8715 3624 8760 3652
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 8938 3652 8944 3664
rect 8812 3624 8944 3652
rect 8812 3612 8818 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 9692 3661 9720 3692
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 10318 3652 10324 3664
rect 9723 3624 10324 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10413 3655 10471 3661
rect 10413 3621 10425 3655
rect 10459 3652 10471 3655
rect 10686 3652 10692 3664
rect 10459 3624 10692 3652
rect 10459 3621 10471 3624
rect 10413 3615 10471 3621
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 4948 3556 5488 3584
rect 5537 3587 5595 3593
rect 4948 3544 4954 3556
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5810 3584 5816 3596
rect 5583 3556 5816 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 9122 3584 9128 3596
rect 7101 3547 7159 3553
rect 7208 3556 9128 3584
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 5626 3516 5632 3528
rect 3099 3488 5632 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 7208 3516 7236 3556
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9824 3587 9882 3593
rect 9824 3553 9836 3587
rect 9870 3584 9882 3587
rect 10594 3584 10600 3596
rect 9870 3556 10600 3584
rect 9870 3553 9882 3556
rect 9824 3547 9882 3553
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 7374 3516 7380 3528
rect 5736 3488 7236 3516
rect 7335 3488 7380 3516
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5736 3448 5764 3488
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 9364 3488 10057 3516
rect 9364 3476 9370 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 5224 3420 5764 3448
rect 5224 3408 5230 3420
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 9953 3451 10011 3457
rect 9953 3448 9965 3451
rect 8168 3420 9965 3448
rect 8168 3408 8174 3420
rect 9953 3417 9965 3420
rect 9999 3417 10011 3451
rect 9953 3411 10011 3417
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 6914 3380 6920 3392
rect 3936 3352 6920 3380
rect 3936 3340 3942 3352
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8128 3380 8156 3408
rect 7524 3352 8156 3380
rect 7524 3340 7530 3352
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 10962 3380 10968 3392
rect 9180 3352 10968 3380
rect 9180 3340 9186 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 1104 3290 11960 3312
rect 1104 3238 2791 3290
rect 2843 3238 2855 3290
rect 2907 3238 2919 3290
rect 2971 3238 2983 3290
rect 3035 3238 6410 3290
rect 6462 3238 6474 3290
rect 6526 3238 6538 3290
rect 6590 3238 6602 3290
rect 6654 3238 10028 3290
rect 10080 3238 10092 3290
rect 10144 3238 10156 3290
rect 10208 3238 10220 3290
rect 10272 3238 11960 3290
rect 1104 3216 11960 3238
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 5258 3176 5264 3188
rect 3559 3148 5264 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 5500 3148 10609 3176
rect 5500 3136 5506 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 5000 3080 7512 3108
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 4890 3040 4896 3052
rect 1995 3012 4896 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 5000 2972 5028 3080
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 7374 3040 7380 3052
rect 5951 3012 7380 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7484 3040 7512 3080
rect 8018 3040 8024 3052
rect 7484 3012 7880 3040
rect 7979 3012 8024 3040
rect 5626 2972 5632 2984
rect 2271 2944 5028 2972
rect 5184 2944 5632 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 5184 2913 5212 2944
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 6880 2944 7757 2972
rect 6880 2932 6886 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7852 2972 7880 3012
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 9398 3040 9404 3052
rect 9359 3012 9404 3040
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9766 2972 9772 2984
rect 7852 2944 9772 2972
rect 7745 2935 7803 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 10318 2972 10324 2984
rect 10279 2944 10324 2972
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 5169 2907 5227 2913
rect 5169 2904 5181 2907
rect 4540 2876 5181 2904
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 4540 2836 4568 2876
rect 5169 2873 5181 2876
rect 5215 2873 5227 2907
rect 5534 2904 5540 2916
rect 5447 2876 5540 2904
rect 5169 2867 5227 2873
rect 5534 2864 5540 2876
rect 5592 2904 5598 2916
rect 7190 2904 7196 2916
rect 5592 2876 7196 2904
rect 5592 2864 5598 2876
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 1820 2808 4568 2836
rect 1820 2796 1826 2808
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 5132 2808 5365 2836
rect 5132 2796 5138 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 7650 2836 7656 2848
rect 5491 2808 7656 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 10520 2836 10548 2935
rect 8076 2808 10548 2836
rect 8076 2796 8082 2808
rect 1104 2746 11960 2768
rect 1104 2694 4600 2746
rect 4652 2694 4664 2746
rect 4716 2694 4728 2746
rect 4780 2694 4792 2746
rect 4844 2694 8219 2746
rect 8271 2694 8283 2746
rect 8335 2694 8347 2746
rect 8399 2694 8411 2746
rect 8463 2694 11960 2746
rect 1104 2672 11960 2694
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 8846 2632 8852 2644
rect 5552 2604 8852 2632
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 3142 2564 3148 2576
rect 2179 2536 3148 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 5552 2564 5580 2604
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 4264 2536 5580 2564
rect 6917 2567 6975 2573
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1544 2499 1602 2505
rect 1544 2465 1556 2499
rect 1590 2496 1602 2499
rect 3878 2496 3884 2508
rect 1590 2468 3884 2496
rect 1590 2465 1602 2468
rect 1544 2459 1602 2465
rect 1412 2360 1440 2459
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4264 2505 4292 2536
rect 6917 2533 6929 2567
rect 6963 2564 6975 2567
rect 7098 2564 7104 2576
rect 6963 2536 7104 2564
rect 6963 2533 6975 2536
rect 6917 2527 6975 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 9769 2567 9827 2573
rect 9769 2533 9781 2567
rect 9815 2564 9827 2567
rect 9858 2564 9864 2576
rect 9815 2536 9864 2564
rect 9815 2533 9827 2536
rect 9769 2527 9827 2533
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 10962 2564 10968 2576
rect 10336 2536 10968 2564
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5442 2496 5448 2508
rect 5040 2468 5448 2496
rect 5040 2456 5046 2468
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 5626 2496 5632 2508
rect 5583 2468 5632 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7340 2468 7389 2496
rect 7340 2456 7346 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7558 2496 7564 2508
rect 7519 2468 7564 2496
rect 7377 2459 7435 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 10336 2505 10364 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 3786 2428 3792 2440
rect 1811 2400 3792 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 7760 2428 7788 2456
rect 5552 2400 7788 2428
rect 5552 2360 5580 2400
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 10459 2431 10517 2437
rect 10459 2428 10471 2431
rect 8996 2400 10471 2428
rect 8996 2388 9002 2400
rect 10459 2397 10471 2400
rect 10505 2397 10517 2431
rect 10459 2391 10517 2397
rect 7466 2360 7472 2372
rect 1412 2332 5580 2360
rect 5644 2332 7472 2360
rect 1673 2295 1731 2301
rect 1673 2261 1685 2295
rect 1719 2292 1731 2295
rect 5644 2292 5672 2332
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 1719 2264 5672 2292
rect 5721 2295 5779 2301
rect 1719 2261 1731 2264
rect 1673 2255 1731 2261
rect 5721 2261 5733 2295
rect 5767 2292 5779 2295
rect 10612 2292 10640 2459
rect 5767 2264 10640 2292
rect 5767 2261 5779 2264
rect 5721 2255 5779 2261
rect 1104 2202 11960 2224
rect 1104 2150 2791 2202
rect 2843 2150 2855 2202
rect 2907 2150 2919 2202
rect 2971 2150 2983 2202
rect 3035 2150 6410 2202
rect 6462 2150 6474 2202
rect 6526 2150 6538 2202
rect 6590 2150 6602 2202
rect 6654 2150 10028 2202
rect 10080 2150 10092 2202
rect 10144 2150 10156 2202
rect 10208 2150 10220 2202
rect 10272 2150 11960 2202
rect 1104 2128 11960 2150
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 10410 2020 10416 2032
rect 4120 1992 10416 2020
rect 4120 1980 4126 1992
rect 10410 1980 10416 1992
rect 10468 1980 10474 2032
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 9582 1952 9588 1964
rect 7892 1924 9588 1952
rect 7892 1912 7898 1924
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
<< via1 >>
rect 2791 13030 2843 13082
rect 2855 13030 2907 13082
rect 2919 13030 2971 13082
rect 2983 13030 3035 13082
rect 6410 13030 6462 13082
rect 6474 13030 6526 13082
rect 6538 13030 6590 13082
rect 6602 13030 6654 13082
rect 10028 13030 10080 13082
rect 10092 13030 10144 13082
rect 10156 13030 10208 13082
rect 10220 13030 10272 13082
rect 9312 12792 9364 12844
rect 3884 12724 3936 12776
rect 4252 12724 4304 12776
rect 5264 12656 5316 12708
rect 4600 12486 4652 12538
rect 4664 12486 4716 12538
rect 4728 12486 4780 12538
rect 4792 12486 4844 12538
rect 8219 12486 8271 12538
rect 8283 12486 8335 12538
rect 8347 12486 8399 12538
rect 8411 12486 8463 12538
rect 3884 12316 3936 12368
rect 4344 12316 4396 12368
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2412 12248 2464 12300
rect 4528 12248 4580 12300
rect 4160 12180 4212 12232
rect 5356 12180 5408 12232
rect 7012 12248 7064 12300
rect 7748 12248 7800 12300
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 9680 12180 9732 12232
rect 2136 12044 2188 12096
rect 6092 12044 6144 12096
rect 2791 11942 2843 11994
rect 2855 11942 2907 11994
rect 2919 11942 2971 11994
rect 2983 11942 3035 11994
rect 6410 11942 6462 11994
rect 6474 11942 6526 11994
rect 6538 11942 6590 11994
rect 6602 11942 6654 11994
rect 10028 11942 10080 11994
rect 10092 11942 10144 11994
rect 10156 11942 10208 11994
rect 10220 11942 10272 11994
rect 10508 11840 10560 11892
rect 3516 11772 3568 11824
rect 4988 11704 5040 11756
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4528 11636 4580 11688
rect 5908 11772 5960 11824
rect 7564 11772 7616 11824
rect 5448 11704 5500 11756
rect 9864 11772 9916 11824
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 6828 11636 6880 11688
rect 7196 11568 7248 11620
rect 7932 11611 7984 11620
rect 5080 11500 5132 11552
rect 5724 11500 5776 11552
rect 7932 11577 7941 11611
rect 7941 11577 7975 11611
rect 7975 11577 7984 11611
rect 7932 11568 7984 11577
rect 9680 11611 9732 11620
rect 9680 11577 9689 11611
rect 9689 11577 9723 11611
rect 9723 11577 9732 11611
rect 9680 11568 9732 11577
rect 10692 11568 10744 11620
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 7748 11500 7800 11509
rect 8024 11500 8076 11552
rect 10876 11500 10928 11552
rect 4600 11398 4652 11450
rect 4664 11398 4716 11450
rect 4728 11398 4780 11450
rect 4792 11398 4844 11450
rect 8219 11398 8271 11450
rect 8283 11398 8335 11450
rect 8347 11398 8399 11450
rect 8411 11398 8463 11450
rect 3792 11296 3844 11348
rect 3976 11296 4028 11348
rect 6184 11296 6236 11348
rect 8576 11296 8628 11348
rect 9312 11296 9364 11348
rect 3332 11160 3384 11212
rect 3608 11160 3660 11212
rect 4988 11160 5040 11212
rect 8024 11160 8076 11212
rect 3240 11092 3292 11144
rect 6276 11092 6328 11144
rect 8116 11092 8168 11144
rect 9128 11092 9180 11144
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 7564 11024 7616 11076
rect 6920 10956 6972 11008
rect 2791 10854 2843 10906
rect 2855 10854 2907 10906
rect 2919 10854 2971 10906
rect 2983 10854 3035 10906
rect 6410 10854 6462 10906
rect 6474 10854 6526 10906
rect 6538 10854 6590 10906
rect 6602 10854 6654 10906
rect 10028 10854 10080 10906
rect 10092 10854 10144 10906
rect 10156 10854 10208 10906
rect 10220 10854 10272 10906
rect 3792 10752 3844 10804
rect 5724 10752 5776 10804
rect 9680 10752 9732 10804
rect 4344 10684 4396 10736
rect 7932 10684 7984 10736
rect 3240 10616 3292 10668
rect 5356 10616 5408 10668
rect 4068 10548 4120 10600
rect 4896 10548 4948 10600
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 6184 10480 6236 10532
rect 6368 10480 6420 10532
rect 5632 10412 5684 10464
rect 6736 10412 6788 10464
rect 9496 10412 9548 10464
rect 4600 10310 4652 10362
rect 4664 10310 4716 10362
rect 4728 10310 4780 10362
rect 4792 10310 4844 10362
rect 8219 10310 8271 10362
rect 8283 10310 8335 10362
rect 8347 10310 8399 10362
rect 8411 10310 8463 10362
rect 3332 10140 3384 10192
rect 1860 10072 1912 10124
rect 3884 10072 3936 10124
rect 5540 10208 5592 10260
rect 7748 10208 7800 10260
rect 5632 10140 5684 10192
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 6000 10072 6052 10124
rect 3148 10004 3200 10056
rect 4252 10004 4304 10056
rect 6092 10004 6144 10056
rect 6368 10072 6420 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 9312 10072 9364 10124
rect 10968 10140 11020 10192
rect 9220 10004 9272 10056
rect 9772 10004 9824 10056
rect 2504 9979 2556 9988
rect 2504 9945 2513 9979
rect 2513 9945 2547 9979
rect 2547 9945 2556 9979
rect 2504 9936 2556 9945
rect 10876 10072 10928 10124
rect 4344 9868 4396 9920
rect 4712 9868 4764 9920
rect 4988 9868 5040 9920
rect 5540 9868 5592 9920
rect 6736 9868 6788 9920
rect 8944 9868 8996 9920
rect 2791 9766 2843 9818
rect 2855 9766 2907 9818
rect 2919 9766 2971 9818
rect 2983 9766 3035 9818
rect 6410 9766 6462 9818
rect 6474 9766 6526 9818
rect 6538 9766 6590 9818
rect 6602 9766 6654 9818
rect 10028 9766 10080 9818
rect 10092 9766 10144 9818
rect 10156 9766 10208 9818
rect 10220 9766 10272 9818
rect 1860 9664 1912 9716
rect 6092 9664 6144 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 10416 9596 10468 9648
rect 5172 9528 5224 9580
rect 6000 9528 6052 9580
rect 9220 9528 9272 9580
rect 3976 9324 4028 9376
rect 5540 9460 5592 9512
rect 5816 9460 5868 9512
rect 6092 9460 6144 9512
rect 6184 9460 6236 9512
rect 8668 9460 8720 9512
rect 9128 9460 9180 9512
rect 4344 9392 4396 9444
rect 6736 9392 6788 9444
rect 7932 9392 7984 9444
rect 9680 9460 9732 9512
rect 10324 9324 10376 9376
rect 10416 9324 10468 9376
rect 4600 9222 4652 9274
rect 4664 9222 4716 9274
rect 4728 9222 4780 9274
rect 4792 9222 4844 9274
rect 8219 9222 8271 9274
rect 8283 9222 8335 9274
rect 8347 9222 8399 9274
rect 8411 9222 8463 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 4252 9120 4304 9172
rect 3884 9052 3936 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 2320 8984 2372 9036
rect 5540 8984 5592 9036
rect 7380 8984 7432 9036
rect 10416 8984 10468 9036
rect 3240 8916 3292 8968
rect 3976 8916 4028 8968
rect 6000 8916 6052 8968
rect 9404 8916 9456 8968
rect 2964 8848 3016 8900
rect 2688 8780 2740 8832
rect 4252 8780 4304 8832
rect 4528 8780 4580 8832
rect 7012 8780 7064 8832
rect 7288 8780 7340 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 2791 8678 2843 8730
rect 2855 8678 2907 8730
rect 2919 8678 2971 8730
rect 2983 8678 3035 8730
rect 6410 8678 6462 8730
rect 6474 8678 6526 8730
rect 6538 8678 6590 8730
rect 6602 8678 6654 8730
rect 10028 8678 10080 8730
rect 10092 8678 10144 8730
rect 10156 8678 10208 8730
rect 10220 8678 10272 8730
rect 9128 8576 9180 8628
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 6828 8508 6880 8560
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 3700 8372 3752 8424
rect 4528 8440 4580 8492
rect 5724 8440 5776 8492
rect 7472 8440 7524 8492
rect 8760 8440 8812 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9588 8440 9640 8492
rect 3976 8372 4028 8424
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 6092 8372 6144 8424
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 9128 8372 9180 8424
rect 9864 8372 9916 8424
rect 5172 8236 5224 8288
rect 5448 8236 5500 8288
rect 8576 8236 8628 8288
rect 4600 8134 4652 8186
rect 4664 8134 4716 8186
rect 4728 8134 4780 8186
rect 4792 8134 4844 8186
rect 8219 8134 8271 8186
rect 8283 8134 8335 8186
rect 8347 8134 8399 8186
rect 8411 8134 8463 8186
rect 2504 8032 2556 8084
rect 7656 8032 7708 8084
rect 1860 8007 1912 8016
rect 1860 7973 1869 8007
rect 1869 7973 1903 8007
rect 1903 7973 1912 8007
rect 1860 7964 1912 7973
rect 3608 7964 3660 8016
rect 4620 7964 4672 8016
rect 4896 7964 4948 8016
rect 5080 8007 5132 8016
rect 5080 7973 5089 8007
rect 5089 7973 5123 8007
rect 5123 7973 5132 8007
rect 5080 7964 5132 7973
rect 7012 7964 7064 8016
rect 8208 7964 8260 8016
rect 8760 7964 8812 8016
rect 10324 7964 10376 8016
rect 2044 7896 2096 7948
rect 4252 7896 4304 7948
rect 4528 7896 4580 7948
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 6920 7896 6972 7948
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5448 7828 5500 7880
rect 6276 7828 6328 7880
rect 6828 7828 6880 7880
rect 5080 7760 5132 7812
rect 7656 7760 7708 7812
rect 8024 7760 8076 7812
rect 4160 7692 4212 7744
rect 7288 7692 7340 7744
rect 7748 7692 7800 7744
rect 2791 7590 2843 7642
rect 2855 7590 2907 7642
rect 2919 7590 2971 7642
rect 2983 7590 3035 7642
rect 6410 7590 6462 7642
rect 6474 7590 6526 7642
rect 6538 7590 6590 7642
rect 6602 7590 6654 7642
rect 10028 7590 10080 7642
rect 10092 7590 10144 7642
rect 10156 7590 10208 7642
rect 10220 7590 10272 7642
rect 2136 7488 2188 7540
rect 2596 7488 2648 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 9496 7488 9548 7540
rect 4252 7420 4304 7472
rect 8116 7420 8168 7472
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 3424 7284 3476 7336
rect 5172 7352 5224 7404
rect 5448 7352 5500 7404
rect 5724 7284 5776 7336
rect 7288 7284 7340 7336
rect 7472 7284 7524 7336
rect 9588 7352 9640 7404
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 3240 7216 3292 7268
rect 7196 7216 7248 7268
rect 9312 7284 9364 7336
rect 2504 7148 2556 7200
rect 3516 7148 3568 7200
rect 5448 7148 5500 7200
rect 6276 7148 6328 7200
rect 7380 7148 7432 7200
rect 7472 7148 7524 7200
rect 9496 7216 9548 7268
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 4600 7046 4652 7098
rect 4664 7046 4716 7098
rect 4728 7046 4780 7098
rect 4792 7046 4844 7098
rect 8219 7046 8271 7098
rect 8283 7046 8335 7098
rect 8347 7046 8399 7098
rect 8411 7046 8463 7098
rect 5080 6944 5132 6996
rect 9680 6944 9732 6996
rect 10784 6944 10836 6996
rect 3148 6808 3200 6860
rect 3608 6808 3660 6860
rect 4160 6808 4212 6860
rect 5448 6876 5500 6928
rect 6276 6876 6328 6928
rect 7288 6919 7340 6928
rect 7288 6885 7297 6919
rect 7297 6885 7331 6919
rect 7331 6885 7340 6919
rect 7288 6876 7340 6885
rect 3792 6672 3844 6724
rect 4252 6740 4304 6792
rect 5632 6808 5684 6860
rect 7104 6808 7156 6860
rect 4620 6672 4672 6724
rect 5264 6740 5316 6792
rect 6828 6740 6880 6792
rect 5448 6672 5500 6724
rect 6276 6672 6328 6724
rect 8116 6672 8168 6724
rect 9956 6715 10008 6724
rect 3424 6604 3476 6656
rect 9956 6681 9965 6715
rect 9965 6681 9999 6715
rect 9999 6681 10008 6715
rect 9956 6672 10008 6681
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 9680 6604 9732 6656
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 2791 6502 2843 6554
rect 2855 6502 2907 6554
rect 2919 6502 2971 6554
rect 2983 6502 3035 6554
rect 6410 6502 6462 6554
rect 6474 6502 6526 6554
rect 6538 6502 6590 6554
rect 6602 6502 6654 6554
rect 10028 6502 10080 6554
rect 10092 6502 10144 6554
rect 10156 6502 10208 6554
rect 10220 6502 10272 6554
rect 4896 6400 4948 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 5724 6400 5776 6452
rect 8484 6400 8536 6452
rect 3884 6332 3936 6384
rect 3700 6264 3752 6316
rect 5356 6332 5408 6384
rect 5448 6332 5500 6384
rect 9312 6332 9364 6384
rect 9956 6332 10008 6384
rect 10508 6332 10560 6384
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 5540 6264 5592 6316
rect 6828 6264 6880 6316
rect 7564 6264 7616 6316
rect 7932 6307 7984 6316
rect 4804 6196 4856 6248
rect 5356 6196 5408 6248
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 5816 6128 5868 6180
rect 6276 6128 6328 6180
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 9220 6264 9272 6316
rect 7748 6196 7800 6248
rect 8024 6196 8076 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 7932 6128 7984 6180
rect 2688 6060 2740 6112
rect 3608 6060 3660 6112
rect 3700 6060 3752 6112
rect 7564 6060 7616 6112
rect 10508 6196 10560 6248
rect 4600 5958 4652 6010
rect 4664 5958 4716 6010
rect 4728 5958 4780 6010
rect 4792 5958 4844 6010
rect 8219 5958 8271 6010
rect 8283 5958 8335 6010
rect 8347 5958 8399 6010
rect 8411 5958 8463 6010
rect 3148 5856 3200 5908
rect 3608 5856 3660 5908
rect 4068 5831 4120 5840
rect 4068 5797 4077 5831
rect 4077 5797 4111 5831
rect 4111 5797 4120 5831
rect 4068 5788 4120 5797
rect 4160 5788 4212 5840
rect 2228 5720 2280 5772
rect 3700 5720 3752 5772
rect 4252 5720 4304 5772
rect 4988 5720 5040 5772
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5264 5763 5316 5772
rect 5080 5720 5132 5729
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6184 5720 6236 5772
rect 6552 5720 6604 5772
rect 7472 5788 7524 5840
rect 8208 5788 8260 5840
rect 7932 5720 7984 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8392 5788 8444 5840
rect 8760 5788 8812 5840
rect 10600 5788 10652 5840
rect 8116 5720 8168 5729
rect 9312 5720 9364 5772
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 3148 5652 3200 5704
rect 1400 5584 1452 5636
rect 2412 5584 2464 5636
rect 8668 5652 8720 5704
rect 9220 5652 9272 5704
rect 7288 5584 7340 5636
rect 8116 5584 8168 5636
rect 6828 5516 6880 5568
rect 8024 5516 8076 5568
rect 8576 5516 8628 5568
rect 9496 5516 9548 5568
rect 2791 5414 2843 5466
rect 2855 5414 2907 5466
rect 2919 5414 2971 5466
rect 2983 5414 3035 5466
rect 6410 5414 6462 5466
rect 6474 5414 6526 5466
rect 6538 5414 6590 5466
rect 6602 5414 6654 5466
rect 10028 5414 10080 5466
rect 10092 5414 10144 5466
rect 10156 5414 10208 5466
rect 10220 5414 10272 5466
rect 1676 5287 1728 5296
rect 1676 5253 1685 5287
rect 1685 5253 1719 5287
rect 1719 5253 1728 5287
rect 1676 5244 1728 5253
rect 3884 5312 3936 5364
rect 7196 5312 7248 5364
rect 9588 5312 9640 5364
rect 5724 5244 5776 5296
rect 6276 5244 6328 5296
rect 6920 5244 6972 5296
rect 9128 5244 9180 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 3792 5176 3844 5228
rect 9680 5176 9732 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 3332 5108 3384 5160
rect 5172 5108 5224 5160
rect 6644 5108 6696 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 6828 5040 6880 5092
rect 8668 5108 8720 5160
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 9588 5040 9640 5092
rect 10876 5040 10928 5092
rect 9220 4972 9272 5024
rect 4600 4870 4652 4922
rect 4664 4870 4716 4922
rect 4728 4870 4780 4922
rect 4792 4870 4844 4922
rect 8219 4870 8271 4922
rect 8283 4870 8335 4922
rect 8347 4870 8399 4922
rect 8411 4870 8463 4922
rect 1768 4768 1820 4820
rect 1676 4700 1728 4752
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 4160 4700 4212 4752
rect 6276 4768 6328 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 10600 4768 10652 4820
rect 3608 4632 3660 4684
rect 3792 4632 3844 4684
rect 4896 4632 4948 4684
rect 5540 4564 5592 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 9772 4700 9824 4752
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 7748 4632 7800 4684
rect 8208 4675 8260 4684
rect 8208 4641 8217 4675
rect 8217 4641 8251 4675
rect 8251 4641 8260 4675
rect 8208 4632 8260 4641
rect 6184 4564 6236 4616
rect 7932 4564 7984 4616
rect 9496 4632 9548 4684
rect 10324 4632 10376 4684
rect 4988 4496 5040 4548
rect 3976 4428 4028 4480
rect 5264 4428 5316 4480
rect 9036 4496 9088 4548
rect 7748 4428 7800 4480
rect 8668 4428 8720 4480
rect 9588 4428 9640 4480
rect 9772 4428 9824 4480
rect 2791 4326 2843 4378
rect 2855 4326 2907 4378
rect 2919 4326 2971 4378
rect 2983 4326 3035 4378
rect 6410 4326 6462 4378
rect 6474 4326 6526 4378
rect 6538 4326 6590 4378
rect 6602 4326 6654 4378
rect 10028 4326 10080 4378
rect 10092 4326 10144 4378
rect 10156 4326 10208 4378
rect 10220 4326 10272 4378
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2596 4156 2648 4208
rect 7012 4224 7064 4276
rect 9496 4224 9548 4276
rect 3424 4088 3476 4140
rect 6184 4156 6236 4208
rect 7932 4156 7984 4208
rect 8208 4156 8260 4208
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 6736 4088 6788 4140
rect 7196 4088 7248 4140
rect 9220 4156 9272 4208
rect 8852 4088 8904 4140
rect 9588 4088 9640 4140
rect 2320 4020 2372 4072
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 5724 4020 5776 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7380 4020 7432 4072
rect 8944 4020 8996 4072
rect 10784 3952 10836 4004
rect 5632 3884 5684 3936
rect 4600 3782 4652 3834
rect 4664 3782 4716 3834
rect 4728 3782 4780 3834
rect 4792 3782 4844 3834
rect 8219 3782 8271 3834
rect 8283 3782 8335 3834
rect 8347 3782 8399 3834
rect 8411 3782 8463 3834
rect 4252 3680 4304 3732
rect 5080 3680 5132 3732
rect 5540 3680 5592 3732
rect 2320 3612 2372 3664
rect 5356 3655 5408 3664
rect 5356 3621 5365 3655
rect 5365 3621 5399 3655
rect 5399 3621 5408 3655
rect 5356 3612 5408 3621
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 3516 3544 3568 3596
rect 4896 3544 4948 3596
rect 5724 3612 5776 3664
rect 6092 3612 6144 3664
rect 8760 3655 8812 3664
rect 8760 3621 8769 3655
rect 8769 3621 8803 3655
rect 8803 3621 8812 3655
rect 8760 3612 8812 3621
rect 8944 3612 8996 3664
rect 10324 3612 10376 3664
rect 10692 3612 10744 3664
rect 5816 3544 5868 3596
rect 6828 3544 6880 3596
rect 5632 3476 5684 3528
rect 9128 3544 9180 3596
rect 10600 3544 10652 3596
rect 7380 3519 7432 3528
rect 5172 3408 5224 3460
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 9312 3476 9364 3528
rect 8116 3408 8168 3460
rect 3884 3340 3936 3392
rect 6920 3340 6972 3392
rect 7472 3340 7524 3392
rect 9128 3340 9180 3392
rect 10968 3340 11020 3392
rect 2791 3238 2843 3290
rect 2855 3238 2907 3290
rect 2919 3238 2971 3290
rect 2983 3238 3035 3290
rect 6410 3238 6462 3290
rect 6474 3238 6526 3290
rect 6538 3238 6590 3290
rect 6602 3238 6654 3290
rect 10028 3238 10080 3290
rect 10092 3238 10144 3290
rect 10156 3238 10208 3290
rect 10220 3238 10272 3290
rect 5264 3136 5316 3188
rect 5448 3136 5500 3188
rect 4896 3000 4948 3052
rect 7380 3000 7432 3052
rect 8024 3043 8076 3052
rect 5632 2932 5684 2984
rect 6828 2932 6880 2984
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 9772 2932 9824 2984
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 1768 2796 1820 2848
rect 5540 2907 5592 2916
rect 5540 2873 5549 2907
rect 5549 2873 5583 2907
rect 5583 2873 5592 2907
rect 5540 2864 5592 2873
rect 7196 2864 7248 2916
rect 5080 2796 5132 2848
rect 7656 2796 7708 2848
rect 8024 2796 8076 2848
rect 4600 2694 4652 2746
rect 4664 2694 4716 2746
rect 4728 2694 4780 2746
rect 4792 2694 4844 2746
rect 8219 2694 8271 2746
rect 8283 2694 8335 2746
rect 8347 2694 8399 2746
rect 8411 2694 8463 2746
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 3148 2524 3200 2576
rect 8852 2592 8904 2644
rect 3884 2456 3936 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 7104 2524 7156 2576
rect 9864 2524 9916 2576
rect 4988 2456 5040 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 5632 2456 5684 2508
rect 7288 2456 7340 2508
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 10968 2524 11020 2576
rect 3792 2388 3844 2440
rect 8944 2388 8996 2440
rect 7472 2320 7524 2372
rect 2791 2150 2843 2202
rect 2855 2150 2907 2202
rect 2919 2150 2971 2202
rect 2983 2150 3035 2202
rect 6410 2150 6462 2202
rect 6474 2150 6526 2202
rect 6538 2150 6590 2202
rect 6602 2150 6654 2202
rect 10028 2150 10080 2202
rect 10092 2150 10144 2202
rect 10156 2150 10208 2202
rect 10220 2150 10272 2202
rect 4068 1980 4120 2032
rect 10416 1980 10468 2032
rect 7840 1912 7892 1964
rect 9588 1912 9640 1964
<< metal2 >>
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 8850 13696 8906 13705
rect 8850 13631 8906 13640
rect 2765 13084 3061 13104
rect 2821 13082 2845 13084
rect 2901 13082 2925 13084
rect 2981 13082 3005 13084
rect 2843 13030 2845 13082
rect 2907 13030 2919 13082
rect 2981 13030 2983 13082
rect 2821 13028 2845 13030
rect 2901 13028 2925 13030
rect 2981 13028 3005 13030
rect 2765 13008 3061 13028
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1412 8430 1440 10639
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 9722 1900 10066
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1674 9480 1730 9489
rect 1674 9415 1730 9424
rect 1688 9042 1716 9415
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1412 5166 1440 5578
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1596 4570 1624 8502
rect 1872 8022 1900 9658
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 2056 7954 2084 10950
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2148 7546 2176 12038
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2240 5778 2268 12242
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 7585 2360 8978
rect 2318 7576 2374 7585
rect 2318 7511 2374 7520
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2240 5658 2268 5714
rect 2240 5630 2360 5658
rect 2424 5642 2452 12242
rect 2765 11996 3061 12016
rect 2821 11994 2845 11996
rect 2901 11994 2925 11996
rect 2981 11994 3005 11996
rect 2843 11942 2845 11994
rect 2907 11942 2919 11994
rect 2981 11942 2983 11994
rect 2821 11940 2845 11942
rect 2901 11940 2925 11942
rect 2981 11940 3005 11942
rect 2765 11920 3061 11940
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2765 10908 3061 10928
rect 2821 10906 2845 10908
rect 2901 10906 2925 10908
rect 2981 10906 3005 10908
rect 2843 10854 2845 10906
rect 2907 10854 2919 10906
rect 2981 10854 2983 10906
rect 2821 10852 2845 10854
rect 2901 10852 2925 10854
rect 2981 10852 3005 10854
rect 2765 10832 3061 10852
rect 3252 10674 3280 11086
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 8090 2544 9930
rect 2765 9820 3061 9840
rect 2821 9818 2845 9820
rect 2901 9818 2925 9820
rect 2981 9818 3005 9820
rect 2843 9766 2845 9818
rect 2907 9766 2919 9818
rect 2981 9766 2983 9818
rect 2821 9764 2845 9766
rect 2901 9764 2925 9766
rect 2981 9764 3005 9766
rect 2765 9744 3061 9764
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2976 8906 3004 9114
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2516 7206 2544 8026
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1688 4758 1716 5238
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1780 4826 1808 5170
rect 2136 5160 2188 5166
rect 2134 5128 2136 5137
rect 2188 5128 2190 5137
rect 2134 5063 2190 5072
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 2332 4690 2360 5630
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1596 4542 1808 4570
rect 1780 3602 1808 4542
rect 2332 4078 2360 4626
rect 2608 4214 2636 7482
rect 2700 6118 2728 8774
rect 2765 8732 3061 8752
rect 2821 8730 2845 8732
rect 2901 8730 2925 8732
rect 2981 8730 3005 8732
rect 2843 8678 2845 8730
rect 2907 8678 2919 8730
rect 2981 8678 2983 8730
rect 2821 8676 2845 8678
rect 2901 8676 2925 8678
rect 2981 8676 3005 8678
rect 2765 8656 3061 8676
rect 2765 7644 3061 7664
rect 2821 7642 2845 7644
rect 2901 7642 2925 7644
rect 2981 7642 3005 7644
rect 2843 7590 2845 7642
rect 2907 7590 2919 7642
rect 2981 7590 2983 7642
rect 2821 7588 2845 7590
rect 2901 7588 2925 7590
rect 2981 7588 3005 7590
rect 2765 7568 3061 7588
rect 3160 7342 3188 9998
rect 3252 8974 3280 10610
rect 3344 10198 3372 11154
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2765 6556 3061 6576
rect 2821 6554 2845 6556
rect 2901 6554 2925 6556
rect 2981 6554 3005 6556
rect 2843 6502 2845 6554
rect 2907 6502 2919 6554
rect 2981 6502 2983 6554
rect 2821 6500 2845 6502
rect 2901 6500 2925 6502
rect 2981 6500 3005 6502
rect 2765 6480 3061 6500
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 3160 5914 3188 6802
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2765 5468 3061 5488
rect 2821 5466 2845 5468
rect 2901 5466 2925 5468
rect 2981 5466 3005 5468
rect 2843 5414 2845 5466
rect 2907 5414 2919 5466
rect 2981 5414 2983 5466
rect 2821 5412 2845 5414
rect 2901 5412 2925 5414
rect 2981 5412 3005 5414
rect 2765 5392 3061 5412
rect 2765 4380 3061 4400
rect 2821 4378 2845 4380
rect 2901 4378 2925 4380
rect 2981 4378 3005 4380
rect 2843 4326 2845 4378
rect 2907 4326 2919 4378
rect 2981 4326 2983 4378
rect 2821 4324 2845 4326
rect 2901 4324 2925 4326
rect 2981 4324 3005 4326
rect 2765 4304 3061 4324
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 1952 4072 2004 4078
rect 1950 4040 1952 4049
rect 2320 4072 2372 4078
rect 2004 4040 2006 4049
rect 2320 4014 2372 4020
rect 1950 3975 2006 3984
rect 2332 3670 2360 4014
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 2854 1808 3538
rect 2765 3292 3061 3312
rect 2821 3290 2845 3292
rect 2901 3290 2925 3292
rect 2981 3290 3005 3292
rect 2843 3238 2845 3290
rect 2907 3238 2919 3290
rect 2981 3238 2983 3290
rect 2821 3236 2845 3238
rect 2901 3236 2925 3238
rect 2981 3236 3005 3238
rect 2765 3216 3061 3236
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 3160 2582 3188 5646
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 2765 2204 3061 2224
rect 2821 2202 2845 2204
rect 2901 2202 2925 2204
rect 2981 2202 3005 2204
rect 2843 2150 2845 2202
rect 2907 2150 2919 2202
rect 2981 2150 2983 2202
rect 2821 2148 2845 2150
rect 2901 2148 2925 2150
rect 2981 2148 3005 2150
rect 2765 2128 3061 2148
rect 3252 200 3280 7210
rect 3344 5166 3372 10134
rect 3436 9761 3464 13631
rect 6384 13084 6680 13104
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6462 13030 6464 13082
rect 6526 13030 6538 13082
rect 6600 13030 6602 13082
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6384 13008 6680 13028
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 3896 12374 3924 12718
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3422 9752 3478 9761
rect 3422 9687 3478 9696
rect 3528 7834 3556 11766
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11354 4016 11630
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3620 8022 3648 11154
rect 3804 10810 3832 11290
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3528 7806 3648 7834
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 6662 3464 7278
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3436 4146 3464 6598
rect 3528 4593 3556 7142
rect 3620 6866 3648 7806
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3712 6322 3740 8366
rect 3804 6882 3832 10746
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 9110 3924 10066
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3988 8974 4016 9318
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3804 6854 3924 6882
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3700 6112 3752 6118
rect 3804 6100 3832 6666
rect 3896 6390 3924 6854
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3752 6072 3832 6100
rect 3700 6054 3752 6060
rect 3620 5914 3648 6054
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3620 4690 3648 5850
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3514 4584 3570 4593
rect 3514 4519 3570 4528
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3528 3602 3556 4519
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3712 1601 3740 5714
rect 3804 5234 3832 6072
rect 3896 5370 3924 6190
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 2446 3832 4626
rect 3988 4486 4016 8366
rect 4080 5846 4108 10542
rect 4172 7886 4200 12174
rect 4264 10062 4292 12718
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 4574 12540 4870 12560
rect 4630 12538 4654 12540
rect 4710 12538 4734 12540
rect 4790 12538 4814 12540
rect 4652 12486 4654 12538
rect 4716 12486 4728 12538
rect 4790 12486 4792 12538
rect 4630 12484 4654 12486
rect 4710 12484 4734 12486
rect 4790 12484 4814 12486
rect 4574 12464 4870 12484
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4356 10742 4384 12310
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4540 11694 4568 12242
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4574 11452 4870 11472
rect 4630 11450 4654 11452
rect 4710 11450 4734 11452
rect 4790 11450 4814 11452
rect 4652 11398 4654 11450
rect 4716 11398 4728 11450
rect 4790 11398 4792 11450
rect 4630 11396 4654 11398
rect 4710 11396 4734 11398
rect 4790 11396 4814 11398
rect 4574 11376 4870 11396
rect 5000 11218 5028 11698
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4264 9178 4292 9998
rect 4356 9926 4384 10678
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4574 10364 4870 10384
rect 4630 10362 4654 10364
rect 4710 10362 4734 10364
rect 4790 10362 4814 10364
rect 4652 10310 4654 10362
rect 4716 10310 4728 10362
rect 4790 10310 4792 10362
rect 4630 10308 4654 10310
rect 4710 10308 4734 10310
rect 4790 10308 4814 10310
rect 4574 10288 4870 10308
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9625 4752 9862
rect 4710 9616 4766 9625
rect 4710 9551 4766 9560
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8537 4292 8774
rect 4250 8528 4306 8537
rect 4250 8463 4306 8472
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 6866 4200 7686
rect 4264 7478 4292 7890
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4172 4758 4200 5782
rect 4264 5778 4292 6734
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4250 5672 4306 5681
rect 4250 5607 4306 5616
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 4264 3738 4292 5607
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 2514 3924 3334
rect 4356 2650 4384 9386
rect 4574 9276 4870 9296
rect 4630 9274 4654 9276
rect 4710 9274 4734 9276
rect 4790 9274 4814 9276
rect 4652 9222 4654 9274
rect 4716 9222 4728 9274
rect 4790 9222 4792 9274
rect 4630 9220 4654 9222
rect 4710 9220 4734 9222
rect 4790 9220 4814 9222
rect 4574 9200 4870 9220
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8498 4568 8774
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4574 8188 4870 8208
rect 4630 8186 4654 8188
rect 4710 8186 4734 8188
rect 4790 8186 4814 8188
rect 4652 8134 4654 8186
rect 4716 8134 4728 8186
rect 4790 8134 4792 8186
rect 4630 8132 4654 8134
rect 4710 8132 4734 8134
rect 4790 8132 4814 8134
rect 4574 8112 4870 8132
rect 4908 8022 4936 10542
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4620 8016 4672 8022
rect 4618 7984 4620 7993
rect 4896 8016 4948 8022
rect 4672 7984 4674 7993
rect 4528 7948 4580 7954
rect 4896 7958 4948 7964
rect 4618 7919 4674 7928
rect 4528 7890 4580 7896
rect 4540 7857 4568 7890
rect 4896 7880 4948 7886
rect 4526 7848 4582 7857
rect 4896 7822 4948 7828
rect 4526 7783 4582 7792
rect 4574 7100 4870 7120
rect 4630 7098 4654 7100
rect 4710 7098 4734 7100
rect 4790 7098 4814 7100
rect 4652 7046 4654 7098
rect 4716 7046 4728 7098
rect 4790 7046 4792 7098
rect 4630 7044 4654 7046
rect 4710 7044 4734 7046
rect 4790 7044 4814 7046
rect 4574 7024 4870 7044
rect 4618 6896 4674 6905
rect 4618 6831 4674 6840
rect 4632 6730 4660 6831
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4802 6488 4858 6497
rect 4908 6458 4936 7822
rect 4802 6423 4858 6432
rect 4896 6452 4948 6458
rect 4816 6254 4844 6423
rect 4896 6394 4948 6400
rect 4894 6352 4950 6361
rect 4894 6287 4950 6296
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4574 6012 4870 6032
rect 4630 6010 4654 6012
rect 4710 6010 4734 6012
rect 4790 6010 4814 6012
rect 4652 5958 4654 6010
rect 4716 5958 4728 6010
rect 4790 5958 4792 6010
rect 4630 5956 4654 5958
rect 4710 5956 4734 5958
rect 4790 5956 4814 5958
rect 4574 5936 4870 5956
rect 4574 4924 4870 4944
rect 4630 4922 4654 4924
rect 4710 4922 4734 4924
rect 4790 4922 4814 4924
rect 4652 4870 4654 4922
rect 4716 4870 4728 4922
rect 4790 4870 4792 4922
rect 4630 4868 4654 4870
rect 4710 4868 4734 4870
rect 4790 4868 4814 4870
rect 4574 4848 4870 4868
rect 4908 4690 4936 6287
rect 5000 5778 5028 9862
rect 5092 8022 5120 11494
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 8294 5212 9522
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 7002 5120 7754
rect 5184 7410 5212 7890
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5092 5778 5120 6938
rect 5276 6882 5304 12650
rect 8193 12540 8489 12560
rect 8249 12538 8273 12540
rect 8329 12538 8353 12540
rect 8409 12538 8433 12540
rect 8271 12486 8273 12538
rect 8335 12486 8347 12538
rect 8409 12486 8411 12538
rect 8249 12484 8273 12486
rect 8329 12484 8353 12486
rect 8409 12484 8433 12486
rect 8193 12464 8489 12484
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5368 11694 5396 12174
rect 5920 11914 5948 12174
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 5828 11886 5948 11914
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5184 6854 5304 6882
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5184 5166 5212 6854
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 5778 5304 6734
rect 5368 6390 5396 10610
rect 5460 9489 5488 11698
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 10266 5580 11630
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10554 5672 10950
rect 5736 10810 5764 11494
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5644 10526 5764 10554
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10198 5672 10406
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9518 5580 9862
rect 5540 9512 5592 9518
rect 5446 9480 5502 9489
rect 5540 9454 5592 9460
rect 5446 9415 5502 9424
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8424 5500 8430
rect 5446 8392 5448 8401
rect 5500 8392 5502 8401
rect 5446 8327 5502 8336
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 7886 5488 8230
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 7206 5488 7346
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6934 5488 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6390 5488 6666
rect 5552 6458 5580 8978
rect 5644 7041 5672 10134
rect 5736 8616 5764 10526
rect 5828 9518 5856 11886
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5736 8588 5856 8616
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5736 7342 5764 8434
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5630 7032 5686 7041
rect 5630 6967 5686 6976
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5552 6322 5580 6394
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4574 3836 4870 3856
rect 4630 3834 4654 3836
rect 4710 3834 4734 3836
rect 4790 3834 4814 3836
rect 4652 3782 4654 3834
rect 4716 3782 4728 3834
rect 4790 3782 4792 3834
rect 4630 3780 4654 3782
rect 4710 3780 4734 3782
rect 4790 3780 4814 3782
rect 4574 3760 4870 3780
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4908 3058 4936 3538
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4574 2748 4870 2768
rect 4630 2746 4654 2748
rect 4710 2746 4734 2748
rect 4790 2746 4814 2748
rect 4652 2694 4654 2746
rect 4716 2694 4728 2746
rect 4790 2694 4792 2746
rect 4630 2692 4654 2694
rect 4710 2692 4734 2694
rect 4790 2692 4814 2694
rect 4574 2672 4870 2692
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 5000 2514 5028 4490
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5092 2854 5120 3674
rect 5184 3466 5212 4014
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5276 3194 5304 4422
rect 5368 3670 5396 6190
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5460 3194 5488 4014
rect 5552 3738 5580 4558
rect 5644 3942 5672 6802
rect 5736 6458 5764 7278
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6338 5856 8588
rect 5736 6310 5856 6338
rect 5736 5302 5764 6310
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5736 4078 5764 4558
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5644 3534 5672 3878
rect 5736 3670 5764 4014
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5828 3602 5856 6122
rect 5920 4146 5948 11766
rect 6104 10198 6132 12038
rect 6384 11996 6680 12016
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6462 11942 6464 11994
rect 6526 11942 6538 11994
rect 6600 11942 6602 11994
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6384 11920 6680 11940
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6196 10538 6224 11290
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9586 6040 10066
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 9722 6132 9998
rect 6288 9722 6316 11086
rect 6384 10908 6680 10928
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6462 10854 6464 10906
rect 6526 10854 6538 10906
rect 6600 10854 6602 10906
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6384 10832 6680 10852
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6380 10130 6408 10474
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6748 9926 6776 10406
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6384 9820 6680 9840
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6462 9766 6464 9818
rect 6526 9766 6538 9818
rect 6600 9766 6602 9818
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6384 9744 6680 9764
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 4690 6040 8910
rect 6104 8430 6132 9454
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6196 7546 6224 9454
rect 6288 7886 6316 9658
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6384 8732 6680 8752
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6462 8678 6464 8730
rect 6526 8678 6538 8730
rect 6600 8678 6602 8730
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6384 8656 6680 8676
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6384 7644 6680 7664
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6462 7590 6464 7642
rect 6526 7590 6538 7642
rect 6600 7590 6602 7642
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6384 7568 6680 7588
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6090 7032 6146 7041
rect 6090 6967 6146 6976
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6104 3670 6132 6967
rect 6196 5778 6224 7482
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6934 6316 7142
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6288 6186 6316 6666
rect 6384 6556 6680 6576
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6462 6502 6464 6554
rect 6526 6502 6538 6554
rect 6600 6502 6602 6554
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6384 6480 6680 6500
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6184 5772 6236 5778
rect 6552 5772 6604 5778
rect 6184 5714 6236 5720
rect 6288 5732 6552 5760
rect 6288 5302 6316 5732
rect 6552 5714 6604 5720
rect 6384 5468 6680 5488
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6462 5414 6464 5466
rect 6526 5414 6538 5466
rect 6600 5414 6602 5466
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6384 5392 6680 5412
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6642 5264 6698 5273
rect 6288 4826 6316 5238
rect 6642 5199 6698 5208
rect 6656 5166 6684 5199
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 4214 6224 4558
rect 6384 4380 6680 4400
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6462 4326 6464 4378
rect 6526 4326 6538 4378
rect 6600 4326 6602 4378
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6384 4304 6680 4324
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 6748 4146 6776 9386
rect 6840 8566 6868 11630
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6840 7886 6868 8502
rect 6932 7954 6960 10950
rect 7024 8838 7052 12242
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8022 7052 8774
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6322 6868 6734
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5098 6868 5510
rect 6932 5302 6960 7890
rect 7010 7848 7066 7857
rect 7010 7783 7066 7792
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6920 5160 6972 5166
rect 7024 5148 7052 7783
rect 7208 7274 7236 11562
rect 7576 11082 7604 11766
rect 7760 11558 7788 12242
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11370 7788 11494
rect 7668 11342 7788 11370
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 7750 7328 8774
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7342 7328 7686
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7208 6916 7236 7210
rect 7392 7206 7420 8978
rect 7484 8498 7512 10066
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7484 7206 7512 7278
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7288 6928 7340 6934
rect 7208 6888 7288 6916
rect 7288 6870 7340 6876
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6972 5120 7052 5148
rect 6920 5102 6972 5108
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6840 4078 6868 5034
rect 6932 4264 6960 5102
rect 7012 4276 7064 4282
rect 6932 4236 7012 4264
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6840 3602 6868 4014
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 6384 3292 6680 3312
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6462 3238 6464 3290
rect 6526 3238 6538 3290
rect 6600 3238 6602 3290
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6384 3216 6680 3236
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 6840 2990 6868 3538
rect 6932 3398 6960 4236
rect 7012 4218 7064 4224
rect 7116 4049 7144 6802
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7208 4298 7236 5306
rect 7300 4826 7328 5578
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7208 4270 7328 4298
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 5448 2508 5500 2514
rect 5552 2496 5580 2858
rect 5644 2514 5672 2926
rect 7116 2582 7144 3975
rect 7208 2922 7236 4082
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7300 2514 7328 4270
rect 7392 4078 7420 7142
rect 7576 6322 7604 11018
rect 7668 8090 7696 11342
rect 7944 10742 7972 11562
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11218 8064 11494
rect 8193 11452 8489 11472
rect 8249 11450 8273 11452
rect 8329 11450 8353 11452
rect 8409 11450 8433 11452
rect 8271 11398 8273 11450
rect 8335 11398 8347 11450
rect 8409 11398 8411 11450
rect 8249 11396 8273 11398
rect 8329 11396 8353 11398
rect 8409 11396 8433 11398
rect 8193 11376 8489 11396
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5846 7512 6190
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7392 3058 7420 3470
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 5500 2468 5580 2496
rect 5632 2508 5684 2514
rect 5448 2450 5500 2456
rect 5632 2450 5684 2456
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4080 2038 4108 2450
rect 7484 2378 7512 3334
rect 7576 2514 7604 6054
rect 7668 2854 7696 7754
rect 7760 7750 7788 10202
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 6746 7788 7686
rect 7760 6718 7880 6746
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 4690 7788 6190
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7760 2514 7788 4422
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 6384 2204 6680 2224
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6462 2150 6464 2202
rect 6526 2150 6538 2202
rect 6600 2150 6602 2202
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6384 2128 6680 2148
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 7852 1970 7880 6718
rect 7944 6322 7972 9386
rect 8036 8430 8064 11154
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8036 7818 8064 8366
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8128 7478 8156 11086
rect 8193 10364 8489 10384
rect 8249 10362 8273 10364
rect 8329 10362 8353 10364
rect 8409 10362 8433 10364
rect 8271 10310 8273 10362
rect 8335 10310 8347 10362
rect 8409 10310 8411 10362
rect 8249 10308 8273 10310
rect 8329 10308 8353 10310
rect 8409 10308 8433 10310
rect 8193 10288 8489 10308
rect 8193 9276 8489 9296
rect 8249 9274 8273 9276
rect 8329 9274 8353 9276
rect 8409 9274 8433 9276
rect 8271 9222 8273 9274
rect 8335 9222 8347 9274
rect 8409 9222 8411 9274
rect 8249 9220 8273 9222
rect 8329 9220 8353 9222
rect 8409 9220 8433 9222
rect 8193 9200 8489 9220
rect 8588 8378 8616 11290
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8668 9512 8720 9518
rect 8772 9466 8800 10542
rect 8720 9460 8800 9466
rect 8668 9454 8800 9460
rect 8680 9438 8800 9454
rect 8772 8498 8800 9438
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8588 8350 8708 8378
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8193 8188 8489 8208
rect 8249 8186 8273 8188
rect 8329 8186 8353 8188
rect 8409 8186 8433 8188
rect 8271 8134 8273 8186
rect 8335 8134 8347 8186
rect 8409 8134 8411 8186
rect 8249 8132 8273 8134
rect 8329 8132 8353 8134
rect 8409 8132 8433 8134
rect 8193 8112 8489 8132
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8024 7336 8076 7342
rect 8220 7290 8248 7958
rect 8076 7284 8248 7290
rect 8024 7278 8248 7284
rect 8036 7262 8248 7278
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8036 6254 8064 7262
rect 8193 7100 8489 7120
rect 8249 7098 8273 7100
rect 8329 7098 8353 7100
rect 8409 7098 8433 7100
rect 8271 7046 8273 7098
rect 8335 7046 8347 7098
rect 8409 7046 8411 7098
rect 8249 7044 8273 7046
rect 8329 7044 8353 7046
rect 8409 7044 8433 7046
rect 8193 7024 8489 7044
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5778 7972 6122
rect 8128 5778 8156 6666
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6458 8524 6598
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8193 6012 8489 6032
rect 8249 6010 8273 6012
rect 8329 6010 8353 6012
rect 8409 6010 8433 6012
rect 8271 5958 8273 6010
rect 8335 5958 8347 6010
rect 8409 5958 8411 6010
rect 8249 5956 8273 5958
rect 8329 5956 8353 5958
rect 8409 5956 8433 5958
rect 8193 5936 8489 5956
rect 8208 5840 8260 5846
rect 8392 5840 8444 5846
rect 8260 5788 8392 5794
rect 8208 5782 8444 5788
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8116 5772 8168 5778
rect 8220 5766 8432 5782
rect 8116 5714 8168 5720
rect 7944 4622 7972 5714
rect 8128 5642 8156 5714
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 2938 7972 4150
rect 8036 3058 8064 5510
rect 8128 3466 8156 5578
rect 8588 5574 8616 8230
rect 8680 5710 8708 8350
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8772 5846 8800 7958
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8193 4924 8489 4944
rect 8249 4922 8273 4924
rect 8329 4922 8353 4924
rect 8409 4922 8433 4924
rect 8271 4870 8273 4922
rect 8335 4870 8347 4922
rect 8409 4870 8411 4922
rect 8249 4868 8273 4870
rect 8329 4868 8353 4870
rect 8409 4868 8433 4870
rect 8193 4848 8489 4868
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8220 4214 8248 4626
rect 8680 4486 8708 5102
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8193 3836 8489 3856
rect 8249 3834 8273 3836
rect 8329 3834 8353 3836
rect 8409 3834 8433 3836
rect 8271 3782 8273 3834
rect 8335 3782 8347 3834
rect 8409 3782 8411 3834
rect 8249 3780 8273 3782
rect 8329 3780 8353 3782
rect 8409 3780 8433 3782
rect 8193 3760 8489 3780
rect 8772 3670 8800 5782
rect 8864 4146 8892 13631
rect 10002 13084 10298 13104
rect 10058 13082 10082 13084
rect 10138 13082 10162 13084
rect 10218 13082 10242 13084
rect 10080 13030 10082 13082
rect 10144 13030 10156 13082
rect 10218 13030 10220 13082
rect 10058 13028 10082 13030
rect 10138 13028 10162 13030
rect 10218 13028 10242 13030
rect 10002 13008 10298 13028
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9324 11354 9352 12786
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11626 9720 12174
rect 10002 11996 10298 12016
rect 10058 11994 10082 11996
rect 10138 11994 10162 11996
rect 10218 11994 10242 11996
rect 10080 11942 10082 11994
rect 10144 11942 10156 11994
rect 10218 11942 10220 11994
rect 10058 11940 10082 11942
rect 10138 11940 10162 11942
rect 10218 11940 10242 11942
rect 10002 11920 10298 11940
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7944 2910 8064 2938
rect 8036 2854 8064 2910
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8193 2748 8489 2768
rect 8249 2746 8273 2748
rect 8329 2746 8353 2748
rect 8409 2746 8433 2748
rect 8271 2694 8273 2746
rect 8335 2694 8347 2746
rect 8409 2694 8411 2746
rect 8249 2692 8273 2694
rect 8329 2692 8353 2694
rect 8409 2692 8433 2694
rect 8193 2672 8489 2692
rect 8864 2650 8892 4082
rect 8956 4078 8984 9862
rect 9140 9518 9168 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9402 10704 9458 10713
rect 9402 10639 9458 10648
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9586 9260 9998
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 8786 9168 9454
rect 9048 8758 9168 8786
rect 9048 4706 9076 8758
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9140 8430 9168 8570
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 5302 9168 8366
rect 9232 6322 9260 9522
rect 9324 7342 9352 10066
rect 9416 8974 9444 10639
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6390 9352 7278
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9232 5030 9260 5646
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9048 4678 9168 4706
rect 9034 4584 9090 4593
rect 9034 4519 9036 4528
rect 9088 4519 9090 4528
rect 9036 4490 9088 4496
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8956 2446 8984 3606
rect 9140 3602 9168 4678
rect 9232 4214 9260 4966
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9140 3398 9168 3538
rect 9324 3534 9352 5714
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9416 3058 9444 8910
rect 9508 8498 9536 10406
rect 9692 9518 9720 10746
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9508 7274 9536 7482
rect 9600 7449 9628 8434
rect 9586 7440 9642 7449
rect 9586 7375 9588 7384
rect 9640 7375 9642 7384
rect 9588 7346 9640 7352
rect 9600 7315 9628 7346
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 7002 9720 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9508 4690 9536 5510
rect 9600 5370 9628 6190
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9586 5264 9642 5273
rect 9692 5234 9720 6598
rect 9586 5199 9642 5208
rect 9680 5228 9732 5234
rect 9600 5098 9628 5199
rect 9680 5170 9732 5176
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9784 4758 9812 9998
rect 9876 8430 9904 11766
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10002 10908 10298 10928
rect 10058 10906 10082 10908
rect 10138 10906 10162 10908
rect 10218 10906 10242 10908
rect 10080 10854 10082 10906
rect 10144 10854 10156 10906
rect 10218 10854 10220 10906
rect 10058 10852 10082 10854
rect 10138 10852 10162 10854
rect 10218 10852 10242 10854
rect 10002 10832 10298 10852
rect 10002 9820 10298 9840
rect 10058 9818 10082 9820
rect 10138 9818 10162 9820
rect 10218 9818 10242 9820
rect 10080 9766 10082 9818
rect 10144 9766 10156 9818
rect 10218 9766 10220 9818
rect 10058 9764 10082 9766
rect 10138 9764 10162 9766
rect 10218 9764 10242 9766
rect 10002 9744 10298 9764
rect 10428 9654 10456 11086
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10002 8732 10298 8752
rect 10058 8730 10082 8732
rect 10138 8730 10162 8732
rect 10218 8730 10242 8732
rect 10080 8678 10082 8730
rect 10144 8678 10156 8730
rect 10218 8678 10220 8730
rect 10058 8676 10082 8678
rect 10138 8676 10162 8678
rect 10218 8676 10242 8678
rect 10002 8656 10298 8676
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 10336 8022 10364 9318
rect 10428 9042 10456 9318
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10002 7644 10298 7664
rect 10058 7642 10082 7644
rect 10138 7642 10162 7644
rect 10218 7642 10242 7644
rect 10080 7590 10082 7642
rect 10144 7590 10156 7642
rect 10218 7590 10220 7642
rect 10058 7588 10082 7590
rect 10138 7588 10162 7590
rect 10218 7588 10242 7590
rect 10002 7568 10298 7588
rect 9876 6730 9996 6746
rect 9876 6724 10008 6730
rect 9876 6718 9956 6724
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9508 4026 9536 4218
rect 9600 4146 9628 4422
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9508 3998 9720 4026
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9692 2802 9720 3998
rect 9784 2990 9812 4422
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9692 2774 9812 2802
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9600 1601 9628 1906
rect 3698 1592 3754 1601
rect 3698 1527 3754 1536
rect 9586 1592 9642 1601
rect 9586 1527 9642 1536
rect 9784 200 9812 2774
rect 9876 2582 9904 6718
rect 9956 6666 10008 6672
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10002 6556 10298 6576
rect 10058 6554 10082 6556
rect 10138 6554 10162 6556
rect 10218 6554 10242 6556
rect 10080 6502 10082 6554
rect 10144 6502 10156 6554
rect 10218 6502 10220 6554
rect 10058 6500 10082 6502
rect 10138 6500 10162 6502
rect 10218 6500 10242 6502
rect 10002 6480 10298 6500
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9968 5778 9996 6326
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10002 5468 10298 5488
rect 10058 5466 10082 5468
rect 10138 5466 10162 5468
rect 10218 5466 10242 5468
rect 10080 5414 10082 5466
rect 10144 5414 10156 5466
rect 10218 5414 10220 5466
rect 10058 5412 10082 5414
rect 10138 5412 10162 5414
rect 10218 5412 10242 5414
rect 10002 5392 10298 5412
rect 10336 4690 10364 6598
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10002 4380 10298 4400
rect 10058 4378 10082 4380
rect 10138 4378 10162 4380
rect 10218 4378 10242 4380
rect 10080 4326 10082 4378
rect 10144 4326 10156 4378
rect 10218 4326 10220 4378
rect 10058 4324 10082 4326
rect 10138 4324 10162 4326
rect 10218 4324 10242 4326
rect 10002 4304 10298 4324
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10002 3292 10298 3312
rect 10058 3290 10082 3292
rect 10138 3290 10162 3292
rect 10218 3290 10242 3292
rect 10080 3238 10082 3290
rect 10144 3238 10156 3290
rect 10218 3238 10220 3290
rect 10058 3236 10082 3238
rect 10138 3236 10162 3238
rect 10218 3236 10242 3238
rect 10002 3216 10298 3236
rect 10336 2990 10364 3606
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10002 2204 10298 2224
rect 10058 2202 10082 2204
rect 10138 2202 10162 2204
rect 10218 2202 10242 2204
rect 10080 2150 10082 2202
rect 10144 2150 10156 2202
rect 10218 2150 10220 2202
rect 10058 2148 10082 2150
rect 10138 2148 10162 2150
rect 10218 2148 10242 2150
rect 10002 2128 10298 2148
rect 10428 2038 10456 8978
rect 10520 6390 10548 11834
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5137 10548 6190
rect 10612 5846 10640 8774
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10600 5160 10652 5166
rect 10506 5128 10562 5137
rect 10600 5102 10652 5108
rect 10506 5063 10562 5072
rect 10612 4826 10640 5102
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10612 3602 10640 4762
rect 10704 3670 10732 11562
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 10130 10916 11494
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10796 4010 10824 6938
rect 10888 5098 10916 10066
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10980 4593 11008 10134
rect 10966 4584 11022 4593
rect 10966 4519 11022 4528
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10980 2582 11008 3334
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 3238 0 3294 200
rect 9770 0 9826 200
<< via2 >>
rect 3422 13640 3478 13696
rect 8850 13640 8906 13696
rect 2765 13082 2821 13084
rect 2845 13082 2901 13084
rect 2925 13082 2981 13084
rect 3005 13082 3061 13084
rect 2765 13030 2791 13082
rect 2791 13030 2821 13082
rect 2845 13030 2855 13082
rect 2855 13030 2901 13082
rect 2925 13030 2971 13082
rect 2971 13030 2981 13082
rect 3005 13030 3035 13082
rect 3035 13030 3061 13082
rect 2765 13028 2821 13030
rect 2845 13028 2901 13030
rect 2925 13028 2981 13030
rect 3005 13028 3061 13030
rect 1398 10648 1454 10704
rect 1674 9424 1730 9480
rect 2318 7520 2374 7576
rect 2765 11994 2821 11996
rect 2845 11994 2901 11996
rect 2925 11994 2981 11996
rect 3005 11994 3061 11996
rect 2765 11942 2791 11994
rect 2791 11942 2821 11994
rect 2845 11942 2855 11994
rect 2855 11942 2901 11994
rect 2925 11942 2971 11994
rect 2971 11942 2981 11994
rect 3005 11942 3035 11994
rect 3035 11942 3061 11994
rect 2765 11940 2821 11942
rect 2845 11940 2901 11942
rect 2925 11940 2981 11942
rect 3005 11940 3061 11942
rect 2765 10906 2821 10908
rect 2845 10906 2901 10908
rect 2925 10906 2981 10908
rect 3005 10906 3061 10908
rect 2765 10854 2791 10906
rect 2791 10854 2821 10906
rect 2845 10854 2855 10906
rect 2855 10854 2901 10906
rect 2925 10854 2971 10906
rect 2971 10854 2981 10906
rect 3005 10854 3035 10906
rect 3035 10854 3061 10906
rect 2765 10852 2821 10854
rect 2845 10852 2901 10854
rect 2925 10852 2981 10854
rect 3005 10852 3061 10854
rect 2765 9818 2821 9820
rect 2845 9818 2901 9820
rect 2925 9818 2981 9820
rect 3005 9818 3061 9820
rect 2765 9766 2791 9818
rect 2791 9766 2821 9818
rect 2845 9766 2855 9818
rect 2855 9766 2901 9818
rect 2925 9766 2971 9818
rect 2971 9766 2981 9818
rect 3005 9766 3035 9818
rect 3035 9766 3061 9818
rect 2765 9764 2821 9766
rect 2845 9764 2901 9766
rect 2925 9764 2981 9766
rect 3005 9764 3061 9766
rect 2134 5108 2136 5128
rect 2136 5108 2188 5128
rect 2188 5108 2190 5128
rect 2134 5072 2190 5108
rect 2765 8730 2821 8732
rect 2845 8730 2901 8732
rect 2925 8730 2981 8732
rect 3005 8730 3061 8732
rect 2765 8678 2791 8730
rect 2791 8678 2821 8730
rect 2845 8678 2855 8730
rect 2855 8678 2901 8730
rect 2925 8678 2971 8730
rect 2971 8678 2981 8730
rect 3005 8678 3035 8730
rect 3035 8678 3061 8730
rect 2765 8676 2821 8678
rect 2845 8676 2901 8678
rect 2925 8676 2981 8678
rect 3005 8676 3061 8678
rect 2765 7642 2821 7644
rect 2845 7642 2901 7644
rect 2925 7642 2981 7644
rect 3005 7642 3061 7644
rect 2765 7590 2791 7642
rect 2791 7590 2821 7642
rect 2845 7590 2855 7642
rect 2855 7590 2901 7642
rect 2925 7590 2971 7642
rect 2971 7590 2981 7642
rect 3005 7590 3035 7642
rect 3035 7590 3061 7642
rect 2765 7588 2821 7590
rect 2845 7588 2901 7590
rect 2925 7588 2981 7590
rect 3005 7588 3061 7590
rect 2765 6554 2821 6556
rect 2845 6554 2901 6556
rect 2925 6554 2981 6556
rect 3005 6554 3061 6556
rect 2765 6502 2791 6554
rect 2791 6502 2821 6554
rect 2845 6502 2855 6554
rect 2855 6502 2901 6554
rect 2925 6502 2971 6554
rect 2971 6502 2981 6554
rect 3005 6502 3035 6554
rect 3035 6502 3061 6554
rect 2765 6500 2821 6502
rect 2845 6500 2901 6502
rect 2925 6500 2981 6502
rect 3005 6500 3061 6502
rect 2765 5466 2821 5468
rect 2845 5466 2901 5468
rect 2925 5466 2981 5468
rect 3005 5466 3061 5468
rect 2765 5414 2791 5466
rect 2791 5414 2821 5466
rect 2845 5414 2855 5466
rect 2855 5414 2901 5466
rect 2925 5414 2971 5466
rect 2971 5414 2981 5466
rect 3005 5414 3035 5466
rect 3035 5414 3061 5466
rect 2765 5412 2821 5414
rect 2845 5412 2901 5414
rect 2925 5412 2981 5414
rect 3005 5412 3061 5414
rect 2765 4378 2821 4380
rect 2845 4378 2901 4380
rect 2925 4378 2981 4380
rect 3005 4378 3061 4380
rect 2765 4326 2791 4378
rect 2791 4326 2821 4378
rect 2845 4326 2855 4378
rect 2855 4326 2901 4378
rect 2925 4326 2971 4378
rect 2971 4326 2981 4378
rect 3005 4326 3035 4378
rect 3035 4326 3061 4378
rect 2765 4324 2821 4326
rect 2845 4324 2901 4326
rect 2925 4324 2981 4326
rect 3005 4324 3061 4326
rect 1950 4020 1952 4040
rect 1952 4020 2004 4040
rect 2004 4020 2006 4040
rect 1950 3984 2006 4020
rect 2765 3290 2821 3292
rect 2845 3290 2901 3292
rect 2925 3290 2981 3292
rect 3005 3290 3061 3292
rect 2765 3238 2791 3290
rect 2791 3238 2821 3290
rect 2845 3238 2855 3290
rect 2855 3238 2901 3290
rect 2925 3238 2971 3290
rect 2971 3238 2981 3290
rect 3005 3238 3035 3290
rect 3035 3238 3061 3290
rect 2765 3236 2821 3238
rect 2845 3236 2901 3238
rect 2925 3236 2981 3238
rect 3005 3236 3061 3238
rect 2765 2202 2821 2204
rect 2845 2202 2901 2204
rect 2925 2202 2981 2204
rect 3005 2202 3061 2204
rect 2765 2150 2791 2202
rect 2791 2150 2821 2202
rect 2845 2150 2855 2202
rect 2855 2150 2901 2202
rect 2925 2150 2971 2202
rect 2971 2150 2981 2202
rect 3005 2150 3035 2202
rect 3035 2150 3061 2202
rect 2765 2148 2821 2150
rect 2845 2148 2901 2150
rect 2925 2148 2981 2150
rect 3005 2148 3061 2150
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6410 13082
rect 6410 13030 6440 13082
rect 6464 13030 6474 13082
rect 6474 13030 6520 13082
rect 6544 13030 6590 13082
rect 6590 13030 6600 13082
rect 6624 13030 6654 13082
rect 6654 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 3422 9696 3478 9752
rect 3514 4528 3570 4584
rect 4574 12538 4630 12540
rect 4654 12538 4710 12540
rect 4734 12538 4790 12540
rect 4814 12538 4870 12540
rect 4574 12486 4600 12538
rect 4600 12486 4630 12538
rect 4654 12486 4664 12538
rect 4664 12486 4710 12538
rect 4734 12486 4780 12538
rect 4780 12486 4790 12538
rect 4814 12486 4844 12538
rect 4844 12486 4870 12538
rect 4574 12484 4630 12486
rect 4654 12484 4710 12486
rect 4734 12484 4790 12486
rect 4814 12484 4870 12486
rect 4574 11450 4630 11452
rect 4654 11450 4710 11452
rect 4734 11450 4790 11452
rect 4814 11450 4870 11452
rect 4574 11398 4600 11450
rect 4600 11398 4630 11450
rect 4654 11398 4664 11450
rect 4664 11398 4710 11450
rect 4734 11398 4780 11450
rect 4780 11398 4790 11450
rect 4814 11398 4844 11450
rect 4844 11398 4870 11450
rect 4574 11396 4630 11398
rect 4654 11396 4710 11398
rect 4734 11396 4790 11398
rect 4814 11396 4870 11398
rect 4574 10362 4630 10364
rect 4654 10362 4710 10364
rect 4734 10362 4790 10364
rect 4814 10362 4870 10364
rect 4574 10310 4600 10362
rect 4600 10310 4630 10362
rect 4654 10310 4664 10362
rect 4664 10310 4710 10362
rect 4734 10310 4780 10362
rect 4780 10310 4790 10362
rect 4814 10310 4844 10362
rect 4844 10310 4870 10362
rect 4574 10308 4630 10310
rect 4654 10308 4710 10310
rect 4734 10308 4790 10310
rect 4814 10308 4870 10310
rect 4710 9560 4766 9616
rect 4250 8472 4306 8528
rect 4250 5616 4306 5672
rect 4574 9274 4630 9276
rect 4654 9274 4710 9276
rect 4734 9274 4790 9276
rect 4814 9274 4870 9276
rect 4574 9222 4600 9274
rect 4600 9222 4630 9274
rect 4654 9222 4664 9274
rect 4664 9222 4710 9274
rect 4734 9222 4780 9274
rect 4780 9222 4790 9274
rect 4814 9222 4844 9274
rect 4844 9222 4870 9274
rect 4574 9220 4630 9222
rect 4654 9220 4710 9222
rect 4734 9220 4790 9222
rect 4814 9220 4870 9222
rect 4574 8186 4630 8188
rect 4654 8186 4710 8188
rect 4734 8186 4790 8188
rect 4814 8186 4870 8188
rect 4574 8134 4600 8186
rect 4600 8134 4630 8186
rect 4654 8134 4664 8186
rect 4664 8134 4710 8186
rect 4734 8134 4780 8186
rect 4780 8134 4790 8186
rect 4814 8134 4844 8186
rect 4844 8134 4870 8186
rect 4574 8132 4630 8134
rect 4654 8132 4710 8134
rect 4734 8132 4790 8134
rect 4814 8132 4870 8134
rect 4618 7964 4620 7984
rect 4620 7964 4672 7984
rect 4672 7964 4674 7984
rect 4618 7928 4674 7964
rect 4526 7792 4582 7848
rect 4574 7098 4630 7100
rect 4654 7098 4710 7100
rect 4734 7098 4790 7100
rect 4814 7098 4870 7100
rect 4574 7046 4600 7098
rect 4600 7046 4630 7098
rect 4654 7046 4664 7098
rect 4664 7046 4710 7098
rect 4734 7046 4780 7098
rect 4780 7046 4790 7098
rect 4814 7046 4844 7098
rect 4844 7046 4870 7098
rect 4574 7044 4630 7046
rect 4654 7044 4710 7046
rect 4734 7044 4790 7046
rect 4814 7044 4870 7046
rect 4618 6840 4674 6896
rect 4802 6432 4858 6488
rect 4894 6296 4950 6352
rect 4574 6010 4630 6012
rect 4654 6010 4710 6012
rect 4734 6010 4790 6012
rect 4814 6010 4870 6012
rect 4574 5958 4600 6010
rect 4600 5958 4630 6010
rect 4654 5958 4664 6010
rect 4664 5958 4710 6010
rect 4734 5958 4780 6010
rect 4780 5958 4790 6010
rect 4814 5958 4844 6010
rect 4844 5958 4870 6010
rect 4574 5956 4630 5958
rect 4654 5956 4710 5958
rect 4734 5956 4790 5958
rect 4814 5956 4870 5958
rect 4574 4922 4630 4924
rect 4654 4922 4710 4924
rect 4734 4922 4790 4924
rect 4814 4922 4870 4924
rect 4574 4870 4600 4922
rect 4600 4870 4630 4922
rect 4654 4870 4664 4922
rect 4664 4870 4710 4922
rect 4734 4870 4780 4922
rect 4780 4870 4790 4922
rect 4814 4870 4844 4922
rect 4844 4870 4870 4922
rect 4574 4868 4630 4870
rect 4654 4868 4710 4870
rect 4734 4868 4790 4870
rect 4814 4868 4870 4870
rect 8193 12538 8249 12540
rect 8273 12538 8329 12540
rect 8353 12538 8409 12540
rect 8433 12538 8489 12540
rect 8193 12486 8219 12538
rect 8219 12486 8249 12538
rect 8273 12486 8283 12538
rect 8283 12486 8329 12538
rect 8353 12486 8399 12538
rect 8399 12486 8409 12538
rect 8433 12486 8463 12538
rect 8463 12486 8489 12538
rect 8193 12484 8249 12486
rect 8273 12484 8329 12486
rect 8353 12484 8409 12486
rect 8433 12484 8489 12486
rect 5446 9424 5502 9480
rect 5446 8372 5448 8392
rect 5448 8372 5500 8392
rect 5500 8372 5502 8392
rect 5446 8336 5502 8372
rect 5630 6976 5686 7032
rect 4574 3834 4630 3836
rect 4654 3834 4710 3836
rect 4734 3834 4790 3836
rect 4814 3834 4870 3836
rect 4574 3782 4600 3834
rect 4600 3782 4630 3834
rect 4654 3782 4664 3834
rect 4664 3782 4710 3834
rect 4734 3782 4780 3834
rect 4780 3782 4790 3834
rect 4814 3782 4844 3834
rect 4844 3782 4870 3834
rect 4574 3780 4630 3782
rect 4654 3780 4710 3782
rect 4734 3780 4790 3782
rect 4814 3780 4870 3782
rect 4574 2746 4630 2748
rect 4654 2746 4710 2748
rect 4734 2746 4790 2748
rect 4814 2746 4870 2748
rect 4574 2694 4600 2746
rect 4600 2694 4630 2746
rect 4654 2694 4664 2746
rect 4664 2694 4710 2746
rect 4734 2694 4780 2746
rect 4780 2694 4790 2746
rect 4814 2694 4844 2746
rect 4844 2694 4870 2746
rect 4574 2692 4630 2694
rect 4654 2692 4710 2694
rect 4734 2692 4790 2694
rect 4814 2692 4870 2694
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6410 11994
rect 6410 11942 6440 11994
rect 6464 11942 6474 11994
rect 6474 11942 6520 11994
rect 6544 11942 6590 11994
rect 6590 11942 6600 11994
rect 6624 11942 6654 11994
rect 6654 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6410 10906
rect 6410 10854 6440 10906
rect 6464 10854 6474 10906
rect 6474 10854 6520 10906
rect 6544 10854 6590 10906
rect 6590 10854 6600 10906
rect 6624 10854 6654 10906
rect 6654 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6410 9818
rect 6410 9766 6440 9818
rect 6464 9766 6474 9818
rect 6474 9766 6520 9818
rect 6544 9766 6590 9818
rect 6590 9766 6600 9818
rect 6624 9766 6654 9818
rect 6654 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6410 8730
rect 6410 8678 6440 8730
rect 6464 8678 6474 8730
rect 6474 8678 6520 8730
rect 6544 8678 6590 8730
rect 6590 8678 6600 8730
rect 6624 8678 6654 8730
rect 6654 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6410 7642
rect 6410 7590 6440 7642
rect 6464 7590 6474 7642
rect 6474 7590 6520 7642
rect 6544 7590 6590 7642
rect 6590 7590 6600 7642
rect 6624 7590 6654 7642
rect 6654 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 6090 6976 6146 7032
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6410 6554
rect 6410 6502 6440 6554
rect 6464 6502 6474 6554
rect 6474 6502 6520 6554
rect 6544 6502 6590 6554
rect 6590 6502 6600 6554
rect 6624 6502 6654 6554
rect 6654 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6410 5466
rect 6410 5414 6440 5466
rect 6464 5414 6474 5466
rect 6474 5414 6520 5466
rect 6544 5414 6590 5466
rect 6590 5414 6600 5466
rect 6624 5414 6654 5466
rect 6654 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 6642 5208 6698 5264
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6410 4378
rect 6410 4326 6440 4378
rect 6464 4326 6474 4378
rect 6474 4326 6520 4378
rect 6544 4326 6590 4378
rect 6590 4326 6600 4378
rect 6624 4326 6654 4378
rect 6654 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 7010 7792 7066 7848
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6410 3290
rect 6410 3238 6440 3290
rect 6464 3238 6474 3290
rect 6474 3238 6520 3290
rect 6544 3238 6590 3290
rect 6590 3238 6600 3290
rect 6624 3238 6654 3290
rect 6654 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 7102 3984 7158 4040
rect 8193 11450 8249 11452
rect 8273 11450 8329 11452
rect 8353 11450 8409 11452
rect 8433 11450 8489 11452
rect 8193 11398 8219 11450
rect 8219 11398 8249 11450
rect 8273 11398 8283 11450
rect 8283 11398 8329 11450
rect 8353 11398 8399 11450
rect 8399 11398 8409 11450
rect 8433 11398 8463 11450
rect 8463 11398 8489 11450
rect 8193 11396 8249 11398
rect 8273 11396 8329 11398
rect 8353 11396 8409 11398
rect 8433 11396 8489 11398
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6410 2202
rect 6410 2150 6440 2202
rect 6464 2150 6474 2202
rect 6474 2150 6520 2202
rect 6544 2150 6590 2202
rect 6590 2150 6600 2202
rect 6624 2150 6654 2202
rect 6654 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 8193 10362 8249 10364
rect 8273 10362 8329 10364
rect 8353 10362 8409 10364
rect 8433 10362 8489 10364
rect 8193 10310 8219 10362
rect 8219 10310 8249 10362
rect 8273 10310 8283 10362
rect 8283 10310 8329 10362
rect 8353 10310 8399 10362
rect 8399 10310 8409 10362
rect 8433 10310 8463 10362
rect 8463 10310 8489 10362
rect 8193 10308 8249 10310
rect 8273 10308 8329 10310
rect 8353 10308 8409 10310
rect 8433 10308 8489 10310
rect 8193 9274 8249 9276
rect 8273 9274 8329 9276
rect 8353 9274 8409 9276
rect 8433 9274 8489 9276
rect 8193 9222 8219 9274
rect 8219 9222 8249 9274
rect 8273 9222 8283 9274
rect 8283 9222 8329 9274
rect 8353 9222 8399 9274
rect 8399 9222 8409 9274
rect 8433 9222 8463 9274
rect 8463 9222 8489 9274
rect 8193 9220 8249 9222
rect 8273 9220 8329 9222
rect 8353 9220 8409 9222
rect 8433 9220 8489 9222
rect 8193 8186 8249 8188
rect 8273 8186 8329 8188
rect 8353 8186 8409 8188
rect 8433 8186 8489 8188
rect 8193 8134 8219 8186
rect 8219 8134 8249 8186
rect 8273 8134 8283 8186
rect 8283 8134 8329 8186
rect 8353 8134 8399 8186
rect 8399 8134 8409 8186
rect 8433 8134 8463 8186
rect 8463 8134 8489 8186
rect 8193 8132 8249 8134
rect 8273 8132 8329 8134
rect 8353 8132 8409 8134
rect 8433 8132 8489 8134
rect 8193 7098 8249 7100
rect 8273 7098 8329 7100
rect 8353 7098 8409 7100
rect 8433 7098 8489 7100
rect 8193 7046 8219 7098
rect 8219 7046 8249 7098
rect 8273 7046 8283 7098
rect 8283 7046 8329 7098
rect 8353 7046 8399 7098
rect 8399 7046 8409 7098
rect 8433 7046 8463 7098
rect 8463 7046 8489 7098
rect 8193 7044 8249 7046
rect 8273 7044 8329 7046
rect 8353 7044 8409 7046
rect 8433 7044 8489 7046
rect 8193 6010 8249 6012
rect 8273 6010 8329 6012
rect 8353 6010 8409 6012
rect 8433 6010 8489 6012
rect 8193 5958 8219 6010
rect 8219 5958 8249 6010
rect 8273 5958 8283 6010
rect 8283 5958 8329 6010
rect 8353 5958 8399 6010
rect 8399 5958 8409 6010
rect 8433 5958 8463 6010
rect 8463 5958 8489 6010
rect 8193 5956 8249 5958
rect 8273 5956 8329 5958
rect 8353 5956 8409 5958
rect 8433 5956 8489 5958
rect 8193 4922 8249 4924
rect 8273 4922 8329 4924
rect 8353 4922 8409 4924
rect 8433 4922 8489 4924
rect 8193 4870 8219 4922
rect 8219 4870 8249 4922
rect 8273 4870 8283 4922
rect 8283 4870 8329 4922
rect 8353 4870 8399 4922
rect 8399 4870 8409 4922
rect 8433 4870 8463 4922
rect 8463 4870 8489 4922
rect 8193 4868 8249 4870
rect 8273 4868 8329 4870
rect 8353 4868 8409 4870
rect 8433 4868 8489 4870
rect 8193 3834 8249 3836
rect 8273 3834 8329 3836
rect 8353 3834 8409 3836
rect 8433 3834 8489 3836
rect 8193 3782 8219 3834
rect 8219 3782 8249 3834
rect 8273 3782 8283 3834
rect 8283 3782 8329 3834
rect 8353 3782 8399 3834
rect 8399 3782 8409 3834
rect 8433 3782 8463 3834
rect 8463 3782 8489 3834
rect 8193 3780 8249 3782
rect 8273 3780 8329 3782
rect 8353 3780 8409 3782
rect 8433 3780 8489 3782
rect 10002 13082 10058 13084
rect 10082 13082 10138 13084
rect 10162 13082 10218 13084
rect 10242 13082 10298 13084
rect 10002 13030 10028 13082
rect 10028 13030 10058 13082
rect 10082 13030 10092 13082
rect 10092 13030 10138 13082
rect 10162 13030 10208 13082
rect 10208 13030 10218 13082
rect 10242 13030 10272 13082
rect 10272 13030 10298 13082
rect 10002 13028 10058 13030
rect 10082 13028 10138 13030
rect 10162 13028 10218 13030
rect 10242 13028 10298 13030
rect 10002 11994 10058 11996
rect 10082 11994 10138 11996
rect 10162 11994 10218 11996
rect 10242 11994 10298 11996
rect 10002 11942 10028 11994
rect 10028 11942 10058 11994
rect 10082 11942 10092 11994
rect 10092 11942 10138 11994
rect 10162 11942 10208 11994
rect 10208 11942 10218 11994
rect 10242 11942 10272 11994
rect 10272 11942 10298 11994
rect 10002 11940 10058 11942
rect 10082 11940 10138 11942
rect 10162 11940 10218 11942
rect 10242 11940 10298 11942
rect 8193 2746 8249 2748
rect 8273 2746 8329 2748
rect 8353 2746 8409 2748
rect 8433 2746 8489 2748
rect 8193 2694 8219 2746
rect 8219 2694 8249 2746
rect 8273 2694 8283 2746
rect 8283 2694 8329 2746
rect 8353 2694 8399 2746
rect 8399 2694 8409 2746
rect 8433 2694 8463 2746
rect 8463 2694 8489 2746
rect 8193 2692 8249 2694
rect 8273 2692 8329 2694
rect 8353 2692 8409 2694
rect 8433 2692 8489 2694
rect 9402 10648 9458 10704
rect 9034 4548 9090 4584
rect 9034 4528 9036 4548
rect 9036 4528 9088 4548
rect 9088 4528 9090 4548
rect 9586 7404 9642 7440
rect 9586 7384 9588 7404
rect 9588 7384 9640 7404
rect 9640 7384 9642 7404
rect 9586 5208 9642 5264
rect 10002 10906 10058 10908
rect 10082 10906 10138 10908
rect 10162 10906 10218 10908
rect 10242 10906 10298 10908
rect 10002 10854 10028 10906
rect 10028 10854 10058 10906
rect 10082 10854 10092 10906
rect 10092 10854 10138 10906
rect 10162 10854 10208 10906
rect 10208 10854 10218 10906
rect 10242 10854 10272 10906
rect 10272 10854 10298 10906
rect 10002 10852 10058 10854
rect 10082 10852 10138 10854
rect 10162 10852 10218 10854
rect 10242 10852 10298 10854
rect 10002 9818 10058 9820
rect 10082 9818 10138 9820
rect 10162 9818 10218 9820
rect 10242 9818 10298 9820
rect 10002 9766 10028 9818
rect 10028 9766 10058 9818
rect 10082 9766 10092 9818
rect 10092 9766 10138 9818
rect 10162 9766 10208 9818
rect 10208 9766 10218 9818
rect 10242 9766 10272 9818
rect 10272 9766 10298 9818
rect 10002 9764 10058 9766
rect 10082 9764 10138 9766
rect 10162 9764 10218 9766
rect 10242 9764 10298 9766
rect 10002 8730 10058 8732
rect 10082 8730 10138 8732
rect 10162 8730 10218 8732
rect 10242 8730 10298 8732
rect 10002 8678 10028 8730
rect 10028 8678 10058 8730
rect 10082 8678 10092 8730
rect 10092 8678 10138 8730
rect 10162 8678 10208 8730
rect 10208 8678 10218 8730
rect 10242 8678 10272 8730
rect 10272 8678 10298 8730
rect 10002 8676 10058 8678
rect 10082 8676 10138 8678
rect 10162 8676 10218 8678
rect 10242 8676 10298 8678
rect 10002 7642 10058 7644
rect 10082 7642 10138 7644
rect 10162 7642 10218 7644
rect 10242 7642 10298 7644
rect 10002 7590 10028 7642
rect 10028 7590 10058 7642
rect 10082 7590 10092 7642
rect 10092 7590 10138 7642
rect 10162 7590 10208 7642
rect 10208 7590 10218 7642
rect 10242 7590 10272 7642
rect 10272 7590 10298 7642
rect 10002 7588 10058 7590
rect 10082 7588 10138 7590
rect 10162 7588 10218 7590
rect 10242 7588 10298 7590
rect 3698 1536 3754 1592
rect 9586 1536 9642 1592
rect 10002 6554 10058 6556
rect 10082 6554 10138 6556
rect 10162 6554 10218 6556
rect 10242 6554 10298 6556
rect 10002 6502 10028 6554
rect 10028 6502 10058 6554
rect 10082 6502 10092 6554
rect 10092 6502 10138 6554
rect 10162 6502 10208 6554
rect 10208 6502 10218 6554
rect 10242 6502 10272 6554
rect 10272 6502 10298 6554
rect 10002 6500 10058 6502
rect 10082 6500 10138 6502
rect 10162 6500 10218 6502
rect 10242 6500 10298 6502
rect 10002 5466 10058 5468
rect 10082 5466 10138 5468
rect 10162 5466 10218 5468
rect 10242 5466 10298 5468
rect 10002 5414 10028 5466
rect 10028 5414 10058 5466
rect 10082 5414 10092 5466
rect 10092 5414 10138 5466
rect 10162 5414 10208 5466
rect 10208 5414 10218 5466
rect 10242 5414 10272 5466
rect 10272 5414 10298 5466
rect 10002 5412 10058 5414
rect 10082 5412 10138 5414
rect 10162 5412 10218 5414
rect 10242 5412 10298 5414
rect 10002 4378 10058 4380
rect 10082 4378 10138 4380
rect 10162 4378 10218 4380
rect 10242 4378 10298 4380
rect 10002 4326 10028 4378
rect 10028 4326 10058 4378
rect 10082 4326 10092 4378
rect 10092 4326 10138 4378
rect 10162 4326 10208 4378
rect 10208 4326 10218 4378
rect 10242 4326 10272 4378
rect 10272 4326 10298 4378
rect 10002 4324 10058 4326
rect 10082 4324 10138 4326
rect 10162 4324 10218 4326
rect 10242 4324 10298 4326
rect 10002 3290 10058 3292
rect 10082 3290 10138 3292
rect 10162 3290 10218 3292
rect 10242 3290 10298 3292
rect 10002 3238 10028 3290
rect 10028 3238 10058 3290
rect 10082 3238 10092 3290
rect 10092 3238 10138 3290
rect 10162 3238 10208 3290
rect 10208 3238 10218 3290
rect 10242 3238 10272 3290
rect 10272 3238 10298 3290
rect 10002 3236 10058 3238
rect 10082 3236 10138 3238
rect 10162 3236 10218 3238
rect 10242 3236 10298 3238
rect 10002 2202 10058 2204
rect 10082 2202 10138 2204
rect 10162 2202 10218 2204
rect 10242 2202 10298 2204
rect 10002 2150 10028 2202
rect 10028 2150 10058 2202
rect 10082 2150 10092 2202
rect 10092 2150 10138 2202
rect 10162 2150 10208 2202
rect 10208 2150 10218 2202
rect 10242 2150 10272 2202
rect 10272 2150 10298 2202
rect 10002 2148 10058 2150
rect 10082 2148 10138 2150
rect 10162 2148 10218 2150
rect 10242 2148 10298 2150
rect 10506 5072 10562 5128
rect 10966 4528 11022 4584
<< metal3 >>
rect 0 13698 200 13728
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13608 200 13638
rect 3417 13635 3483 13638
rect 8845 13698 8911 13701
rect 12902 13698 13102 13728
rect 8845 13696 13102 13698
rect 8845 13640 8850 13696
rect 8906 13640 13102 13696
rect 8845 13638 13102 13640
rect 8845 13635 8911 13638
rect 12902 13608 13102 13638
rect 2753 13088 3073 13089
rect 2753 13024 2761 13088
rect 2825 13024 2841 13088
rect 2905 13024 2921 13088
rect 2985 13024 3001 13088
rect 3065 13024 3073 13088
rect 2753 13023 3073 13024
rect 6372 13088 6692 13089
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 13023 6692 13024
rect 9990 13088 10310 13089
rect 9990 13024 9998 13088
rect 10062 13024 10078 13088
rect 10142 13024 10158 13088
rect 10222 13024 10238 13088
rect 10302 13024 10310 13088
rect 9990 13023 10310 13024
rect 4562 12544 4882 12545
rect 4562 12480 4570 12544
rect 4634 12480 4650 12544
rect 4714 12480 4730 12544
rect 4794 12480 4810 12544
rect 4874 12480 4882 12544
rect 4562 12479 4882 12480
rect 8181 12544 8501 12545
rect 8181 12480 8189 12544
rect 8253 12480 8269 12544
rect 8333 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8501 12544
rect 8181 12479 8501 12480
rect 2753 12000 3073 12001
rect 2753 11936 2761 12000
rect 2825 11936 2841 12000
rect 2905 11936 2921 12000
rect 2985 11936 3001 12000
rect 3065 11936 3073 12000
rect 2753 11935 3073 11936
rect 6372 12000 6692 12001
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 11935 6692 11936
rect 9990 12000 10310 12001
rect 9990 11936 9998 12000
rect 10062 11936 10078 12000
rect 10142 11936 10158 12000
rect 10222 11936 10238 12000
rect 10302 11936 10310 12000
rect 9990 11935 10310 11936
rect 4562 11456 4882 11457
rect 4562 11392 4570 11456
rect 4634 11392 4650 11456
rect 4714 11392 4730 11456
rect 4794 11392 4810 11456
rect 4874 11392 4882 11456
rect 4562 11391 4882 11392
rect 8181 11456 8501 11457
rect 8181 11392 8189 11456
rect 8253 11392 8269 11456
rect 8333 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8501 11456
rect 8181 11391 8501 11392
rect 2753 10912 3073 10913
rect 2753 10848 2761 10912
rect 2825 10848 2841 10912
rect 2905 10848 2921 10912
rect 2985 10848 3001 10912
rect 3065 10848 3073 10912
rect 2753 10847 3073 10848
rect 6372 10912 6692 10913
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 10847 6692 10848
rect 9990 10912 10310 10913
rect 9990 10848 9998 10912
rect 10062 10848 10078 10912
rect 10142 10848 10158 10912
rect 10222 10848 10238 10912
rect 10302 10848 10310 10912
rect 9990 10847 10310 10848
rect 0 10706 200 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 200 10646
rect 1393 10643 1459 10646
rect 9397 10706 9463 10709
rect 12902 10706 13102 10736
rect 9397 10704 13102 10706
rect 9397 10648 9402 10704
rect 9458 10648 13102 10704
rect 9397 10646 13102 10648
rect 9397 10643 9463 10646
rect 12902 10616 13102 10646
rect 4562 10368 4882 10369
rect 4562 10304 4570 10368
rect 4634 10304 4650 10368
rect 4714 10304 4730 10368
rect 4794 10304 4810 10368
rect 4874 10304 4882 10368
rect 4562 10303 4882 10304
rect 8181 10368 8501 10369
rect 8181 10304 8189 10368
rect 8253 10304 8269 10368
rect 8333 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8501 10368
rect 8181 10303 8501 10304
rect 2753 9824 3073 9825
rect 2753 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2921 9824
rect 2985 9760 3001 9824
rect 3065 9760 3073 9824
rect 2753 9759 3073 9760
rect 6372 9824 6692 9825
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 9759 6692 9760
rect 9990 9824 10310 9825
rect 9990 9760 9998 9824
rect 10062 9760 10078 9824
rect 10142 9760 10158 9824
rect 10222 9760 10238 9824
rect 10302 9760 10310 9824
rect 9990 9759 10310 9760
rect 3417 9754 3483 9757
rect 3417 9752 4538 9754
rect 3417 9696 3422 9752
rect 3478 9696 4538 9752
rect 3417 9694 4538 9696
rect 3417 9691 3483 9694
rect 4102 9556 4108 9620
rect 4172 9618 4178 9620
rect 4478 9618 4538 9694
rect 4172 9558 4538 9618
rect 4705 9618 4771 9621
rect 5022 9618 5028 9620
rect 4705 9616 5028 9618
rect 4705 9560 4710 9616
rect 4766 9560 5028 9616
rect 4705 9558 5028 9560
rect 4172 9556 4178 9558
rect 4705 9555 4771 9558
rect 5022 9556 5028 9558
rect 5092 9556 5098 9620
rect 1669 9482 1735 9485
rect 5441 9482 5507 9485
rect 1669 9480 5507 9482
rect 1669 9424 1674 9480
rect 1730 9424 5446 9480
rect 5502 9424 5507 9480
rect 1669 9422 5507 9424
rect 1669 9419 1735 9422
rect 5441 9419 5507 9422
rect 4562 9280 4882 9281
rect 4562 9216 4570 9280
rect 4634 9216 4650 9280
rect 4714 9216 4730 9280
rect 4794 9216 4810 9280
rect 4874 9216 4882 9280
rect 4562 9215 4882 9216
rect 8181 9280 8501 9281
rect 8181 9216 8189 9280
rect 8253 9216 8269 9280
rect 8333 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8501 9280
rect 8181 9215 8501 9216
rect 2753 8736 3073 8737
rect 2753 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2921 8736
rect 2985 8672 3001 8736
rect 3065 8672 3073 8736
rect 2753 8671 3073 8672
rect 6372 8736 6692 8737
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 8671 6692 8672
rect 9990 8736 10310 8737
rect 9990 8672 9998 8736
rect 10062 8672 10078 8736
rect 10142 8672 10158 8736
rect 10222 8672 10238 8736
rect 10302 8672 10310 8736
rect 9990 8671 10310 8672
rect 4245 8532 4311 8533
rect 4245 8530 4292 8532
rect 4200 8528 4292 8530
rect 4200 8472 4250 8528
rect 4200 8470 4292 8472
rect 4245 8468 4292 8470
rect 4356 8468 4362 8532
rect 4245 8467 4311 8468
rect 5441 8394 5507 8397
rect 5398 8392 5507 8394
rect 5398 8336 5446 8392
rect 5502 8336 5507 8392
rect 5398 8331 5507 8336
rect 4562 8192 4882 8193
rect 4562 8128 4570 8192
rect 4634 8128 4650 8192
rect 4714 8128 4730 8192
rect 4794 8128 4810 8192
rect 4874 8128 4882 8192
rect 4562 8127 4882 8128
rect 4286 7924 4292 7988
rect 4356 7986 4362 7988
rect 4613 7986 4679 7989
rect 4356 7984 4679 7986
rect 4356 7928 4618 7984
rect 4674 7928 4679 7984
rect 4356 7926 4679 7928
rect 4356 7924 4362 7926
rect 4613 7923 4679 7926
rect 4521 7850 4587 7853
rect 5398 7850 5458 8331
rect 8181 8192 8501 8193
rect 8181 8128 8189 8192
rect 8253 8128 8269 8192
rect 8333 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8501 8192
rect 8181 8127 8501 8128
rect 7005 7850 7071 7853
rect 4521 7848 7071 7850
rect 4521 7792 4526 7848
rect 4582 7792 7010 7848
rect 7066 7792 7071 7848
rect 4521 7790 7071 7792
rect 4521 7787 4587 7790
rect 7005 7787 7071 7790
rect 2753 7648 3073 7649
rect 0 7578 200 7608
rect 2753 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2921 7648
rect 2985 7584 3001 7648
rect 3065 7584 3073 7648
rect 2753 7583 3073 7584
rect 6372 7648 6692 7649
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 7583 6692 7584
rect 9990 7648 10310 7649
rect 9990 7584 9998 7648
rect 10062 7584 10078 7648
rect 10142 7584 10158 7648
rect 10222 7584 10238 7648
rect 10302 7584 10310 7648
rect 9990 7583 10310 7584
rect 2313 7578 2379 7581
rect 12902 7578 13102 7608
rect 0 7576 2379 7578
rect 0 7520 2318 7576
rect 2374 7520 2379 7576
rect 0 7518 2379 7520
rect 0 7488 200 7518
rect 2313 7515 2379 7518
rect 10550 7518 13102 7578
rect 9581 7442 9647 7445
rect 10550 7442 10610 7518
rect 12902 7488 13102 7518
rect 9581 7440 10610 7442
rect 9581 7384 9586 7440
rect 9642 7384 10610 7440
rect 9581 7382 10610 7384
rect 9581 7379 9647 7382
rect 4562 7104 4882 7105
rect 4562 7040 4570 7104
rect 4634 7040 4650 7104
rect 4714 7040 4730 7104
rect 4794 7040 4810 7104
rect 4874 7040 4882 7104
rect 4562 7039 4882 7040
rect 8181 7104 8501 7105
rect 8181 7040 8189 7104
rect 8253 7040 8269 7104
rect 8333 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8501 7104
rect 8181 7039 8501 7040
rect 5625 7034 5691 7037
rect 6085 7034 6151 7037
rect 5030 7032 6151 7034
rect 5030 6976 5630 7032
rect 5686 6976 6090 7032
rect 6146 6976 6151 7032
rect 5030 6974 6151 6976
rect 4613 6898 4679 6901
rect 5030 6898 5090 6974
rect 5625 6971 5691 6974
rect 6085 6971 6151 6974
rect 4613 6896 5090 6898
rect 4613 6840 4618 6896
rect 4674 6840 5090 6896
rect 4613 6838 5090 6840
rect 4613 6835 4679 6838
rect 2753 6560 3073 6561
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3073 6560
rect 2753 6495 3073 6496
rect 6372 6560 6692 6561
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 6495 6692 6496
rect 9990 6560 10310 6561
rect 9990 6496 9998 6560
rect 10062 6496 10078 6560
rect 10142 6496 10158 6560
rect 10222 6496 10238 6560
rect 10302 6496 10310 6560
rect 9990 6495 10310 6496
rect 4102 6428 4108 6492
rect 4172 6490 4178 6492
rect 4797 6490 4863 6493
rect 4172 6488 4863 6490
rect 4172 6432 4802 6488
rect 4858 6432 4863 6488
rect 4172 6430 4863 6432
rect 4172 6428 4178 6430
rect 4797 6427 4863 6430
rect 4889 6354 4955 6357
rect 5022 6354 5028 6356
rect 4889 6352 5028 6354
rect 4889 6296 4894 6352
rect 4950 6296 5028 6352
rect 4889 6294 5028 6296
rect 4889 6291 4955 6294
rect 5022 6292 5028 6294
rect 5092 6292 5098 6356
rect 4562 6016 4882 6017
rect 4562 5952 4570 6016
rect 4634 5952 4650 6016
rect 4714 5952 4730 6016
rect 4794 5952 4810 6016
rect 4874 5952 4882 6016
rect 4562 5951 4882 5952
rect 8181 6016 8501 6017
rect 8181 5952 8189 6016
rect 8253 5952 8269 6016
rect 8333 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8501 6016
rect 8181 5951 8501 5952
rect 4245 5676 4311 5677
rect 4245 5672 4292 5676
rect 4356 5674 4362 5676
rect 4245 5616 4250 5672
rect 4245 5612 4292 5616
rect 4356 5614 4402 5674
rect 4356 5612 4362 5614
rect 4245 5611 4311 5612
rect 2753 5472 3073 5473
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3073 5472
rect 2753 5407 3073 5408
rect 6372 5472 6692 5473
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 5407 6692 5408
rect 9990 5472 10310 5473
rect 9990 5408 9998 5472
rect 10062 5408 10078 5472
rect 10142 5408 10158 5472
rect 10222 5408 10238 5472
rect 10302 5408 10310 5472
rect 9990 5407 10310 5408
rect 6637 5266 6703 5269
rect 9581 5266 9647 5269
rect 6637 5264 9647 5266
rect 6637 5208 6642 5264
rect 6698 5208 9586 5264
rect 9642 5208 9647 5264
rect 6637 5206 9647 5208
rect 6637 5203 6703 5206
rect 9581 5203 9647 5206
rect 2129 5130 2195 5133
rect 10501 5130 10567 5133
rect 2129 5128 10567 5130
rect 2129 5072 2134 5128
rect 2190 5072 10506 5128
rect 10562 5072 10567 5128
rect 2129 5070 10567 5072
rect 2129 5067 2195 5070
rect 10501 5067 10567 5070
rect 4562 4928 4882 4929
rect 4562 4864 4570 4928
rect 4634 4864 4650 4928
rect 4714 4864 4730 4928
rect 4794 4864 4810 4928
rect 4874 4864 4882 4928
rect 4562 4863 4882 4864
rect 8181 4928 8501 4929
rect 8181 4864 8189 4928
rect 8253 4864 8269 4928
rect 8333 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8501 4928
rect 8181 4863 8501 4864
rect 0 4586 200 4616
rect 3509 4586 3575 4589
rect 0 4584 3575 4586
rect 0 4528 3514 4584
rect 3570 4528 3575 4584
rect 0 4526 3575 4528
rect 0 4496 200 4526
rect 3509 4523 3575 4526
rect 9029 4586 9095 4589
rect 10961 4586 11027 4589
rect 12902 4586 13102 4616
rect 9029 4584 13102 4586
rect 9029 4528 9034 4584
rect 9090 4528 10966 4584
rect 11022 4528 13102 4584
rect 9029 4526 13102 4528
rect 9029 4523 9095 4526
rect 10961 4523 11027 4526
rect 12902 4496 13102 4526
rect 2753 4384 3073 4385
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3073 4384
rect 2753 4319 3073 4320
rect 6372 4384 6692 4385
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 4319 6692 4320
rect 9990 4384 10310 4385
rect 9990 4320 9998 4384
rect 10062 4320 10078 4384
rect 10142 4320 10158 4384
rect 10222 4320 10238 4384
rect 10302 4320 10310 4384
rect 9990 4319 10310 4320
rect 1945 4042 2011 4045
rect 7097 4042 7163 4045
rect 1945 4040 7163 4042
rect 1945 3984 1950 4040
rect 2006 3984 7102 4040
rect 7158 3984 7163 4040
rect 1945 3982 7163 3984
rect 1945 3979 2011 3982
rect 7097 3979 7163 3982
rect 4562 3840 4882 3841
rect 4562 3776 4570 3840
rect 4634 3776 4650 3840
rect 4714 3776 4730 3840
rect 4794 3776 4810 3840
rect 4874 3776 4882 3840
rect 4562 3775 4882 3776
rect 8181 3840 8501 3841
rect 8181 3776 8189 3840
rect 8253 3776 8269 3840
rect 8333 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8501 3840
rect 8181 3775 8501 3776
rect 2753 3296 3073 3297
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3073 3296
rect 2753 3231 3073 3232
rect 6372 3296 6692 3297
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 3231 6692 3232
rect 9990 3296 10310 3297
rect 9990 3232 9998 3296
rect 10062 3232 10078 3296
rect 10142 3232 10158 3296
rect 10222 3232 10238 3296
rect 10302 3232 10310 3296
rect 9990 3231 10310 3232
rect 4562 2752 4882 2753
rect 4562 2688 4570 2752
rect 4634 2688 4650 2752
rect 4714 2688 4730 2752
rect 4794 2688 4810 2752
rect 4874 2688 4882 2752
rect 4562 2687 4882 2688
rect 8181 2752 8501 2753
rect 8181 2688 8189 2752
rect 8253 2688 8269 2752
rect 8333 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8501 2752
rect 8181 2687 8501 2688
rect 2753 2208 3073 2209
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3073 2208
rect 2753 2143 3073 2144
rect 6372 2208 6692 2209
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2143 6692 2144
rect 9990 2208 10310 2209
rect 9990 2144 9998 2208
rect 10062 2144 10078 2208
rect 10142 2144 10158 2208
rect 10222 2144 10238 2208
rect 10302 2144 10310 2208
rect 9990 2143 10310 2144
rect 0 1594 200 1624
rect 3693 1594 3759 1597
rect 0 1592 3759 1594
rect 0 1536 3698 1592
rect 3754 1536 3759 1592
rect 0 1534 3759 1536
rect 0 1504 200 1534
rect 3693 1531 3759 1534
rect 9581 1594 9647 1597
rect 12902 1594 13102 1624
rect 9581 1592 13102 1594
rect 9581 1536 9586 1592
rect 9642 1536 13102 1592
rect 9581 1534 13102 1536
rect 9581 1531 9647 1534
rect 12902 1504 13102 1534
<< via3 >>
rect 2761 13084 2825 13088
rect 2761 13028 2765 13084
rect 2765 13028 2821 13084
rect 2821 13028 2825 13084
rect 2761 13024 2825 13028
rect 2841 13084 2905 13088
rect 2841 13028 2845 13084
rect 2845 13028 2901 13084
rect 2901 13028 2905 13084
rect 2841 13024 2905 13028
rect 2921 13084 2985 13088
rect 2921 13028 2925 13084
rect 2925 13028 2981 13084
rect 2981 13028 2985 13084
rect 2921 13024 2985 13028
rect 3001 13084 3065 13088
rect 3001 13028 3005 13084
rect 3005 13028 3061 13084
rect 3061 13028 3065 13084
rect 3001 13024 3065 13028
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 9998 13084 10062 13088
rect 9998 13028 10002 13084
rect 10002 13028 10058 13084
rect 10058 13028 10062 13084
rect 9998 13024 10062 13028
rect 10078 13084 10142 13088
rect 10078 13028 10082 13084
rect 10082 13028 10138 13084
rect 10138 13028 10142 13084
rect 10078 13024 10142 13028
rect 10158 13084 10222 13088
rect 10158 13028 10162 13084
rect 10162 13028 10218 13084
rect 10218 13028 10222 13084
rect 10158 13024 10222 13028
rect 10238 13084 10302 13088
rect 10238 13028 10242 13084
rect 10242 13028 10298 13084
rect 10298 13028 10302 13084
rect 10238 13024 10302 13028
rect 4570 12540 4634 12544
rect 4570 12484 4574 12540
rect 4574 12484 4630 12540
rect 4630 12484 4634 12540
rect 4570 12480 4634 12484
rect 4650 12540 4714 12544
rect 4650 12484 4654 12540
rect 4654 12484 4710 12540
rect 4710 12484 4714 12540
rect 4650 12480 4714 12484
rect 4730 12540 4794 12544
rect 4730 12484 4734 12540
rect 4734 12484 4790 12540
rect 4790 12484 4794 12540
rect 4730 12480 4794 12484
rect 4810 12540 4874 12544
rect 4810 12484 4814 12540
rect 4814 12484 4870 12540
rect 4870 12484 4874 12540
rect 4810 12480 4874 12484
rect 8189 12540 8253 12544
rect 8189 12484 8193 12540
rect 8193 12484 8249 12540
rect 8249 12484 8253 12540
rect 8189 12480 8253 12484
rect 8269 12540 8333 12544
rect 8269 12484 8273 12540
rect 8273 12484 8329 12540
rect 8329 12484 8333 12540
rect 8269 12480 8333 12484
rect 8349 12540 8413 12544
rect 8349 12484 8353 12540
rect 8353 12484 8409 12540
rect 8409 12484 8413 12540
rect 8349 12480 8413 12484
rect 8429 12540 8493 12544
rect 8429 12484 8433 12540
rect 8433 12484 8489 12540
rect 8489 12484 8493 12540
rect 8429 12480 8493 12484
rect 2761 11996 2825 12000
rect 2761 11940 2765 11996
rect 2765 11940 2821 11996
rect 2821 11940 2825 11996
rect 2761 11936 2825 11940
rect 2841 11996 2905 12000
rect 2841 11940 2845 11996
rect 2845 11940 2901 11996
rect 2901 11940 2905 11996
rect 2841 11936 2905 11940
rect 2921 11996 2985 12000
rect 2921 11940 2925 11996
rect 2925 11940 2981 11996
rect 2981 11940 2985 11996
rect 2921 11936 2985 11940
rect 3001 11996 3065 12000
rect 3001 11940 3005 11996
rect 3005 11940 3061 11996
rect 3061 11940 3065 11996
rect 3001 11936 3065 11940
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 9998 11996 10062 12000
rect 9998 11940 10002 11996
rect 10002 11940 10058 11996
rect 10058 11940 10062 11996
rect 9998 11936 10062 11940
rect 10078 11996 10142 12000
rect 10078 11940 10082 11996
rect 10082 11940 10138 11996
rect 10138 11940 10142 11996
rect 10078 11936 10142 11940
rect 10158 11996 10222 12000
rect 10158 11940 10162 11996
rect 10162 11940 10218 11996
rect 10218 11940 10222 11996
rect 10158 11936 10222 11940
rect 10238 11996 10302 12000
rect 10238 11940 10242 11996
rect 10242 11940 10298 11996
rect 10298 11940 10302 11996
rect 10238 11936 10302 11940
rect 4570 11452 4634 11456
rect 4570 11396 4574 11452
rect 4574 11396 4630 11452
rect 4630 11396 4634 11452
rect 4570 11392 4634 11396
rect 4650 11452 4714 11456
rect 4650 11396 4654 11452
rect 4654 11396 4710 11452
rect 4710 11396 4714 11452
rect 4650 11392 4714 11396
rect 4730 11452 4794 11456
rect 4730 11396 4734 11452
rect 4734 11396 4790 11452
rect 4790 11396 4794 11452
rect 4730 11392 4794 11396
rect 4810 11452 4874 11456
rect 4810 11396 4814 11452
rect 4814 11396 4870 11452
rect 4870 11396 4874 11452
rect 4810 11392 4874 11396
rect 8189 11452 8253 11456
rect 8189 11396 8193 11452
rect 8193 11396 8249 11452
rect 8249 11396 8253 11452
rect 8189 11392 8253 11396
rect 8269 11452 8333 11456
rect 8269 11396 8273 11452
rect 8273 11396 8329 11452
rect 8329 11396 8333 11452
rect 8269 11392 8333 11396
rect 8349 11452 8413 11456
rect 8349 11396 8353 11452
rect 8353 11396 8409 11452
rect 8409 11396 8413 11452
rect 8349 11392 8413 11396
rect 8429 11452 8493 11456
rect 8429 11396 8433 11452
rect 8433 11396 8489 11452
rect 8489 11396 8493 11452
rect 8429 11392 8493 11396
rect 2761 10908 2825 10912
rect 2761 10852 2765 10908
rect 2765 10852 2821 10908
rect 2821 10852 2825 10908
rect 2761 10848 2825 10852
rect 2841 10908 2905 10912
rect 2841 10852 2845 10908
rect 2845 10852 2901 10908
rect 2901 10852 2905 10908
rect 2841 10848 2905 10852
rect 2921 10908 2985 10912
rect 2921 10852 2925 10908
rect 2925 10852 2981 10908
rect 2981 10852 2985 10908
rect 2921 10848 2985 10852
rect 3001 10908 3065 10912
rect 3001 10852 3005 10908
rect 3005 10852 3061 10908
rect 3061 10852 3065 10908
rect 3001 10848 3065 10852
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 9998 10908 10062 10912
rect 9998 10852 10002 10908
rect 10002 10852 10058 10908
rect 10058 10852 10062 10908
rect 9998 10848 10062 10852
rect 10078 10908 10142 10912
rect 10078 10852 10082 10908
rect 10082 10852 10138 10908
rect 10138 10852 10142 10908
rect 10078 10848 10142 10852
rect 10158 10908 10222 10912
rect 10158 10852 10162 10908
rect 10162 10852 10218 10908
rect 10218 10852 10222 10908
rect 10158 10848 10222 10852
rect 10238 10908 10302 10912
rect 10238 10852 10242 10908
rect 10242 10852 10298 10908
rect 10298 10852 10302 10908
rect 10238 10848 10302 10852
rect 4570 10364 4634 10368
rect 4570 10308 4574 10364
rect 4574 10308 4630 10364
rect 4630 10308 4634 10364
rect 4570 10304 4634 10308
rect 4650 10364 4714 10368
rect 4650 10308 4654 10364
rect 4654 10308 4710 10364
rect 4710 10308 4714 10364
rect 4650 10304 4714 10308
rect 4730 10364 4794 10368
rect 4730 10308 4734 10364
rect 4734 10308 4790 10364
rect 4790 10308 4794 10364
rect 4730 10304 4794 10308
rect 4810 10364 4874 10368
rect 4810 10308 4814 10364
rect 4814 10308 4870 10364
rect 4870 10308 4874 10364
rect 4810 10304 4874 10308
rect 8189 10364 8253 10368
rect 8189 10308 8193 10364
rect 8193 10308 8249 10364
rect 8249 10308 8253 10364
rect 8189 10304 8253 10308
rect 8269 10364 8333 10368
rect 8269 10308 8273 10364
rect 8273 10308 8329 10364
rect 8329 10308 8333 10364
rect 8269 10304 8333 10308
rect 8349 10364 8413 10368
rect 8349 10308 8353 10364
rect 8353 10308 8409 10364
rect 8409 10308 8413 10364
rect 8349 10304 8413 10308
rect 8429 10364 8493 10368
rect 8429 10308 8433 10364
rect 8433 10308 8489 10364
rect 8489 10308 8493 10364
rect 8429 10304 8493 10308
rect 2761 9820 2825 9824
rect 2761 9764 2765 9820
rect 2765 9764 2821 9820
rect 2821 9764 2825 9820
rect 2761 9760 2825 9764
rect 2841 9820 2905 9824
rect 2841 9764 2845 9820
rect 2845 9764 2901 9820
rect 2901 9764 2905 9820
rect 2841 9760 2905 9764
rect 2921 9820 2985 9824
rect 2921 9764 2925 9820
rect 2925 9764 2981 9820
rect 2981 9764 2985 9820
rect 2921 9760 2985 9764
rect 3001 9820 3065 9824
rect 3001 9764 3005 9820
rect 3005 9764 3061 9820
rect 3061 9764 3065 9820
rect 3001 9760 3065 9764
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 9998 9820 10062 9824
rect 9998 9764 10002 9820
rect 10002 9764 10058 9820
rect 10058 9764 10062 9820
rect 9998 9760 10062 9764
rect 10078 9820 10142 9824
rect 10078 9764 10082 9820
rect 10082 9764 10138 9820
rect 10138 9764 10142 9820
rect 10078 9760 10142 9764
rect 10158 9820 10222 9824
rect 10158 9764 10162 9820
rect 10162 9764 10218 9820
rect 10218 9764 10222 9820
rect 10158 9760 10222 9764
rect 10238 9820 10302 9824
rect 10238 9764 10242 9820
rect 10242 9764 10298 9820
rect 10298 9764 10302 9820
rect 10238 9760 10302 9764
rect 4108 9556 4172 9620
rect 5028 9556 5092 9620
rect 4570 9276 4634 9280
rect 4570 9220 4574 9276
rect 4574 9220 4630 9276
rect 4630 9220 4634 9276
rect 4570 9216 4634 9220
rect 4650 9276 4714 9280
rect 4650 9220 4654 9276
rect 4654 9220 4710 9276
rect 4710 9220 4714 9276
rect 4650 9216 4714 9220
rect 4730 9276 4794 9280
rect 4730 9220 4734 9276
rect 4734 9220 4790 9276
rect 4790 9220 4794 9276
rect 4730 9216 4794 9220
rect 4810 9276 4874 9280
rect 4810 9220 4814 9276
rect 4814 9220 4870 9276
rect 4870 9220 4874 9276
rect 4810 9216 4874 9220
rect 8189 9276 8253 9280
rect 8189 9220 8193 9276
rect 8193 9220 8249 9276
rect 8249 9220 8253 9276
rect 8189 9216 8253 9220
rect 8269 9276 8333 9280
rect 8269 9220 8273 9276
rect 8273 9220 8329 9276
rect 8329 9220 8333 9276
rect 8269 9216 8333 9220
rect 8349 9276 8413 9280
rect 8349 9220 8353 9276
rect 8353 9220 8409 9276
rect 8409 9220 8413 9276
rect 8349 9216 8413 9220
rect 8429 9276 8493 9280
rect 8429 9220 8433 9276
rect 8433 9220 8489 9276
rect 8489 9220 8493 9276
rect 8429 9216 8493 9220
rect 2761 8732 2825 8736
rect 2761 8676 2765 8732
rect 2765 8676 2821 8732
rect 2821 8676 2825 8732
rect 2761 8672 2825 8676
rect 2841 8732 2905 8736
rect 2841 8676 2845 8732
rect 2845 8676 2901 8732
rect 2901 8676 2905 8732
rect 2841 8672 2905 8676
rect 2921 8732 2985 8736
rect 2921 8676 2925 8732
rect 2925 8676 2981 8732
rect 2981 8676 2985 8732
rect 2921 8672 2985 8676
rect 3001 8732 3065 8736
rect 3001 8676 3005 8732
rect 3005 8676 3061 8732
rect 3061 8676 3065 8732
rect 3001 8672 3065 8676
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 9998 8732 10062 8736
rect 9998 8676 10002 8732
rect 10002 8676 10058 8732
rect 10058 8676 10062 8732
rect 9998 8672 10062 8676
rect 10078 8732 10142 8736
rect 10078 8676 10082 8732
rect 10082 8676 10138 8732
rect 10138 8676 10142 8732
rect 10078 8672 10142 8676
rect 10158 8732 10222 8736
rect 10158 8676 10162 8732
rect 10162 8676 10218 8732
rect 10218 8676 10222 8732
rect 10158 8672 10222 8676
rect 10238 8732 10302 8736
rect 10238 8676 10242 8732
rect 10242 8676 10298 8732
rect 10298 8676 10302 8732
rect 10238 8672 10302 8676
rect 4292 8528 4356 8532
rect 4292 8472 4306 8528
rect 4306 8472 4356 8528
rect 4292 8468 4356 8472
rect 4570 8188 4634 8192
rect 4570 8132 4574 8188
rect 4574 8132 4630 8188
rect 4630 8132 4634 8188
rect 4570 8128 4634 8132
rect 4650 8188 4714 8192
rect 4650 8132 4654 8188
rect 4654 8132 4710 8188
rect 4710 8132 4714 8188
rect 4650 8128 4714 8132
rect 4730 8188 4794 8192
rect 4730 8132 4734 8188
rect 4734 8132 4790 8188
rect 4790 8132 4794 8188
rect 4730 8128 4794 8132
rect 4810 8188 4874 8192
rect 4810 8132 4814 8188
rect 4814 8132 4870 8188
rect 4870 8132 4874 8188
rect 4810 8128 4874 8132
rect 4292 7924 4356 7988
rect 8189 8188 8253 8192
rect 8189 8132 8193 8188
rect 8193 8132 8249 8188
rect 8249 8132 8253 8188
rect 8189 8128 8253 8132
rect 8269 8188 8333 8192
rect 8269 8132 8273 8188
rect 8273 8132 8329 8188
rect 8329 8132 8333 8188
rect 8269 8128 8333 8132
rect 8349 8188 8413 8192
rect 8349 8132 8353 8188
rect 8353 8132 8409 8188
rect 8409 8132 8413 8188
rect 8349 8128 8413 8132
rect 8429 8188 8493 8192
rect 8429 8132 8433 8188
rect 8433 8132 8489 8188
rect 8489 8132 8493 8188
rect 8429 8128 8493 8132
rect 2761 7644 2825 7648
rect 2761 7588 2765 7644
rect 2765 7588 2821 7644
rect 2821 7588 2825 7644
rect 2761 7584 2825 7588
rect 2841 7644 2905 7648
rect 2841 7588 2845 7644
rect 2845 7588 2901 7644
rect 2901 7588 2905 7644
rect 2841 7584 2905 7588
rect 2921 7644 2985 7648
rect 2921 7588 2925 7644
rect 2925 7588 2981 7644
rect 2981 7588 2985 7644
rect 2921 7584 2985 7588
rect 3001 7644 3065 7648
rect 3001 7588 3005 7644
rect 3005 7588 3061 7644
rect 3061 7588 3065 7644
rect 3001 7584 3065 7588
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 9998 7644 10062 7648
rect 9998 7588 10002 7644
rect 10002 7588 10058 7644
rect 10058 7588 10062 7644
rect 9998 7584 10062 7588
rect 10078 7644 10142 7648
rect 10078 7588 10082 7644
rect 10082 7588 10138 7644
rect 10138 7588 10142 7644
rect 10078 7584 10142 7588
rect 10158 7644 10222 7648
rect 10158 7588 10162 7644
rect 10162 7588 10218 7644
rect 10218 7588 10222 7644
rect 10158 7584 10222 7588
rect 10238 7644 10302 7648
rect 10238 7588 10242 7644
rect 10242 7588 10298 7644
rect 10298 7588 10302 7644
rect 10238 7584 10302 7588
rect 4570 7100 4634 7104
rect 4570 7044 4574 7100
rect 4574 7044 4630 7100
rect 4630 7044 4634 7100
rect 4570 7040 4634 7044
rect 4650 7100 4714 7104
rect 4650 7044 4654 7100
rect 4654 7044 4710 7100
rect 4710 7044 4714 7100
rect 4650 7040 4714 7044
rect 4730 7100 4794 7104
rect 4730 7044 4734 7100
rect 4734 7044 4790 7100
rect 4790 7044 4794 7100
rect 4730 7040 4794 7044
rect 4810 7100 4874 7104
rect 4810 7044 4814 7100
rect 4814 7044 4870 7100
rect 4870 7044 4874 7100
rect 4810 7040 4874 7044
rect 8189 7100 8253 7104
rect 8189 7044 8193 7100
rect 8193 7044 8249 7100
rect 8249 7044 8253 7100
rect 8189 7040 8253 7044
rect 8269 7100 8333 7104
rect 8269 7044 8273 7100
rect 8273 7044 8329 7100
rect 8329 7044 8333 7100
rect 8269 7040 8333 7044
rect 8349 7100 8413 7104
rect 8349 7044 8353 7100
rect 8353 7044 8409 7100
rect 8409 7044 8413 7100
rect 8349 7040 8413 7044
rect 8429 7100 8493 7104
rect 8429 7044 8433 7100
rect 8433 7044 8489 7100
rect 8489 7044 8493 7100
rect 8429 7040 8493 7044
rect 2761 6556 2825 6560
rect 2761 6500 2765 6556
rect 2765 6500 2821 6556
rect 2821 6500 2825 6556
rect 2761 6496 2825 6500
rect 2841 6556 2905 6560
rect 2841 6500 2845 6556
rect 2845 6500 2901 6556
rect 2901 6500 2905 6556
rect 2841 6496 2905 6500
rect 2921 6556 2985 6560
rect 2921 6500 2925 6556
rect 2925 6500 2981 6556
rect 2981 6500 2985 6556
rect 2921 6496 2985 6500
rect 3001 6556 3065 6560
rect 3001 6500 3005 6556
rect 3005 6500 3061 6556
rect 3061 6500 3065 6556
rect 3001 6496 3065 6500
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 9998 6556 10062 6560
rect 9998 6500 10002 6556
rect 10002 6500 10058 6556
rect 10058 6500 10062 6556
rect 9998 6496 10062 6500
rect 10078 6556 10142 6560
rect 10078 6500 10082 6556
rect 10082 6500 10138 6556
rect 10138 6500 10142 6556
rect 10078 6496 10142 6500
rect 10158 6556 10222 6560
rect 10158 6500 10162 6556
rect 10162 6500 10218 6556
rect 10218 6500 10222 6556
rect 10158 6496 10222 6500
rect 10238 6556 10302 6560
rect 10238 6500 10242 6556
rect 10242 6500 10298 6556
rect 10298 6500 10302 6556
rect 10238 6496 10302 6500
rect 4108 6428 4172 6492
rect 5028 6292 5092 6356
rect 4570 6012 4634 6016
rect 4570 5956 4574 6012
rect 4574 5956 4630 6012
rect 4630 5956 4634 6012
rect 4570 5952 4634 5956
rect 4650 6012 4714 6016
rect 4650 5956 4654 6012
rect 4654 5956 4710 6012
rect 4710 5956 4714 6012
rect 4650 5952 4714 5956
rect 4730 6012 4794 6016
rect 4730 5956 4734 6012
rect 4734 5956 4790 6012
rect 4790 5956 4794 6012
rect 4730 5952 4794 5956
rect 4810 6012 4874 6016
rect 4810 5956 4814 6012
rect 4814 5956 4870 6012
rect 4870 5956 4874 6012
rect 4810 5952 4874 5956
rect 8189 6012 8253 6016
rect 8189 5956 8193 6012
rect 8193 5956 8249 6012
rect 8249 5956 8253 6012
rect 8189 5952 8253 5956
rect 8269 6012 8333 6016
rect 8269 5956 8273 6012
rect 8273 5956 8329 6012
rect 8329 5956 8333 6012
rect 8269 5952 8333 5956
rect 8349 6012 8413 6016
rect 8349 5956 8353 6012
rect 8353 5956 8409 6012
rect 8409 5956 8413 6012
rect 8349 5952 8413 5956
rect 8429 6012 8493 6016
rect 8429 5956 8433 6012
rect 8433 5956 8489 6012
rect 8489 5956 8493 6012
rect 8429 5952 8493 5956
rect 4292 5672 4356 5676
rect 4292 5616 4306 5672
rect 4306 5616 4356 5672
rect 4292 5612 4356 5616
rect 2761 5468 2825 5472
rect 2761 5412 2765 5468
rect 2765 5412 2821 5468
rect 2821 5412 2825 5468
rect 2761 5408 2825 5412
rect 2841 5468 2905 5472
rect 2841 5412 2845 5468
rect 2845 5412 2901 5468
rect 2901 5412 2905 5468
rect 2841 5408 2905 5412
rect 2921 5468 2985 5472
rect 2921 5412 2925 5468
rect 2925 5412 2981 5468
rect 2981 5412 2985 5468
rect 2921 5408 2985 5412
rect 3001 5468 3065 5472
rect 3001 5412 3005 5468
rect 3005 5412 3061 5468
rect 3061 5412 3065 5468
rect 3001 5408 3065 5412
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 9998 5468 10062 5472
rect 9998 5412 10002 5468
rect 10002 5412 10058 5468
rect 10058 5412 10062 5468
rect 9998 5408 10062 5412
rect 10078 5468 10142 5472
rect 10078 5412 10082 5468
rect 10082 5412 10138 5468
rect 10138 5412 10142 5468
rect 10078 5408 10142 5412
rect 10158 5468 10222 5472
rect 10158 5412 10162 5468
rect 10162 5412 10218 5468
rect 10218 5412 10222 5468
rect 10158 5408 10222 5412
rect 10238 5468 10302 5472
rect 10238 5412 10242 5468
rect 10242 5412 10298 5468
rect 10298 5412 10302 5468
rect 10238 5408 10302 5412
rect 4570 4924 4634 4928
rect 4570 4868 4574 4924
rect 4574 4868 4630 4924
rect 4630 4868 4634 4924
rect 4570 4864 4634 4868
rect 4650 4924 4714 4928
rect 4650 4868 4654 4924
rect 4654 4868 4710 4924
rect 4710 4868 4714 4924
rect 4650 4864 4714 4868
rect 4730 4924 4794 4928
rect 4730 4868 4734 4924
rect 4734 4868 4790 4924
rect 4790 4868 4794 4924
rect 4730 4864 4794 4868
rect 4810 4924 4874 4928
rect 4810 4868 4814 4924
rect 4814 4868 4870 4924
rect 4870 4868 4874 4924
rect 4810 4864 4874 4868
rect 8189 4924 8253 4928
rect 8189 4868 8193 4924
rect 8193 4868 8249 4924
rect 8249 4868 8253 4924
rect 8189 4864 8253 4868
rect 8269 4924 8333 4928
rect 8269 4868 8273 4924
rect 8273 4868 8329 4924
rect 8329 4868 8333 4924
rect 8269 4864 8333 4868
rect 8349 4924 8413 4928
rect 8349 4868 8353 4924
rect 8353 4868 8409 4924
rect 8409 4868 8413 4924
rect 8349 4864 8413 4868
rect 8429 4924 8493 4928
rect 8429 4868 8433 4924
rect 8433 4868 8489 4924
rect 8489 4868 8493 4924
rect 8429 4864 8493 4868
rect 2761 4380 2825 4384
rect 2761 4324 2765 4380
rect 2765 4324 2821 4380
rect 2821 4324 2825 4380
rect 2761 4320 2825 4324
rect 2841 4380 2905 4384
rect 2841 4324 2845 4380
rect 2845 4324 2901 4380
rect 2901 4324 2905 4380
rect 2841 4320 2905 4324
rect 2921 4380 2985 4384
rect 2921 4324 2925 4380
rect 2925 4324 2981 4380
rect 2981 4324 2985 4380
rect 2921 4320 2985 4324
rect 3001 4380 3065 4384
rect 3001 4324 3005 4380
rect 3005 4324 3061 4380
rect 3061 4324 3065 4380
rect 3001 4320 3065 4324
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 9998 4380 10062 4384
rect 9998 4324 10002 4380
rect 10002 4324 10058 4380
rect 10058 4324 10062 4380
rect 9998 4320 10062 4324
rect 10078 4380 10142 4384
rect 10078 4324 10082 4380
rect 10082 4324 10138 4380
rect 10138 4324 10142 4380
rect 10078 4320 10142 4324
rect 10158 4380 10222 4384
rect 10158 4324 10162 4380
rect 10162 4324 10218 4380
rect 10218 4324 10222 4380
rect 10158 4320 10222 4324
rect 10238 4380 10302 4384
rect 10238 4324 10242 4380
rect 10242 4324 10298 4380
rect 10298 4324 10302 4380
rect 10238 4320 10302 4324
rect 4570 3836 4634 3840
rect 4570 3780 4574 3836
rect 4574 3780 4630 3836
rect 4630 3780 4634 3836
rect 4570 3776 4634 3780
rect 4650 3836 4714 3840
rect 4650 3780 4654 3836
rect 4654 3780 4710 3836
rect 4710 3780 4714 3836
rect 4650 3776 4714 3780
rect 4730 3836 4794 3840
rect 4730 3780 4734 3836
rect 4734 3780 4790 3836
rect 4790 3780 4794 3836
rect 4730 3776 4794 3780
rect 4810 3836 4874 3840
rect 4810 3780 4814 3836
rect 4814 3780 4870 3836
rect 4870 3780 4874 3836
rect 4810 3776 4874 3780
rect 8189 3836 8253 3840
rect 8189 3780 8193 3836
rect 8193 3780 8249 3836
rect 8249 3780 8253 3836
rect 8189 3776 8253 3780
rect 8269 3836 8333 3840
rect 8269 3780 8273 3836
rect 8273 3780 8329 3836
rect 8329 3780 8333 3836
rect 8269 3776 8333 3780
rect 8349 3836 8413 3840
rect 8349 3780 8353 3836
rect 8353 3780 8409 3836
rect 8409 3780 8413 3836
rect 8349 3776 8413 3780
rect 8429 3836 8493 3840
rect 8429 3780 8433 3836
rect 8433 3780 8489 3836
rect 8489 3780 8493 3836
rect 8429 3776 8493 3780
rect 2761 3292 2825 3296
rect 2761 3236 2765 3292
rect 2765 3236 2821 3292
rect 2821 3236 2825 3292
rect 2761 3232 2825 3236
rect 2841 3292 2905 3296
rect 2841 3236 2845 3292
rect 2845 3236 2901 3292
rect 2901 3236 2905 3292
rect 2841 3232 2905 3236
rect 2921 3292 2985 3296
rect 2921 3236 2925 3292
rect 2925 3236 2981 3292
rect 2981 3236 2985 3292
rect 2921 3232 2985 3236
rect 3001 3292 3065 3296
rect 3001 3236 3005 3292
rect 3005 3236 3061 3292
rect 3061 3236 3065 3292
rect 3001 3232 3065 3236
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 9998 3292 10062 3296
rect 9998 3236 10002 3292
rect 10002 3236 10058 3292
rect 10058 3236 10062 3292
rect 9998 3232 10062 3236
rect 10078 3292 10142 3296
rect 10078 3236 10082 3292
rect 10082 3236 10138 3292
rect 10138 3236 10142 3292
rect 10078 3232 10142 3236
rect 10158 3292 10222 3296
rect 10158 3236 10162 3292
rect 10162 3236 10218 3292
rect 10218 3236 10222 3292
rect 10158 3232 10222 3236
rect 10238 3292 10302 3296
rect 10238 3236 10242 3292
rect 10242 3236 10298 3292
rect 10298 3236 10302 3292
rect 10238 3232 10302 3236
rect 4570 2748 4634 2752
rect 4570 2692 4574 2748
rect 4574 2692 4630 2748
rect 4630 2692 4634 2748
rect 4570 2688 4634 2692
rect 4650 2748 4714 2752
rect 4650 2692 4654 2748
rect 4654 2692 4710 2748
rect 4710 2692 4714 2748
rect 4650 2688 4714 2692
rect 4730 2748 4794 2752
rect 4730 2692 4734 2748
rect 4734 2692 4790 2748
rect 4790 2692 4794 2748
rect 4730 2688 4794 2692
rect 4810 2748 4874 2752
rect 4810 2692 4814 2748
rect 4814 2692 4870 2748
rect 4870 2692 4874 2748
rect 4810 2688 4874 2692
rect 8189 2748 8253 2752
rect 8189 2692 8193 2748
rect 8193 2692 8249 2748
rect 8249 2692 8253 2748
rect 8189 2688 8253 2692
rect 8269 2748 8333 2752
rect 8269 2692 8273 2748
rect 8273 2692 8329 2748
rect 8329 2692 8333 2748
rect 8269 2688 8333 2692
rect 8349 2748 8413 2752
rect 8349 2692 8353 2748
rect 8353 2692 8409 2748
rect 8409 2692 8413 2748
rect 8349 2688 8413 2692
rect 8429 2748 8493 2752
rect 8429 2692 8433 2748
rect 8433 2692 8489 2748
rect 8489 2692 8493 2748
rect 8429 2688 8493 2692
rect 2761 2204 2825 2208
rect 2761 2148 2765 2204
rect 2765 2148 2821 2204
rect 2821 2148 2825 2204
rect 2761 2144 2825 2148
rect 2841 2204 2905 2208
rect 2841 2148 2845 2204
rect 2845 2148 2901 2204
rect 2901 2148 2905 2204
rect 2841 2144 2905 2148
rect 2921 2204 2985 2208
rect 2921 2148 2925 2204
rect 2925 2148 2981 2204
rect 2981 2148 2985 2204
rect 2921 2144 2985 2148
rect 3001 2204 3065 2208
rect 3001 2148 3005 2204
rect 3005 2148 3061 2204
rect 3061 2148 3065 2204
rect 3001 2144 3065 2148
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 9998 2204 10062 2208
rect 9998 2148 10002 2204
rect 10002 2148 10058 2204
rect 10058 2148 10062 2204
rect 9998 2144 10062 2148
rect 10078 2204 10142 2208
rect 10078 2148 10082 2204
rect 10082 2148 10138 2204
rect 10138 2148 10142 2204
rect 10078 2144 10142 2148
rect 10158 2204 10222 2208
rect 10158 2148 10162 2204
rect 10162 2148 10218 2204
rect 10218 2148 10222 2204
rect 10158 2144 10222 2148
rect 10238 2204 10302 2208
rect 10238 2148 10242 2204
rect 10242 2148 10298 2204
rect 10298 2148 10302 2204
rect 10238 2144 10302 2148
<< metal4 >>
rect 2753 13088 3073 13104
rect 2753 13024 2761 13088
rect 2825 13024 2841 13088
rect 2905 13024 2921 13088
rect 2985 13024 3001 13088
rect 3065 13024 3073 13088
rect 2753 12000 3073 13024
rect 2753 11936 2761 12000
rect 2825 11936 2841 12000
rect 2905 11936 2921 12000
rect 2985 11936 3001 12000
rect 3065 11936 3073 12000
rect 2753 11312 3073 11936
rect 2753 11076 2795 11312
rect 3031 11076 3073 11312
rect 2753 10912 3073 11076
rect 2753 10848 2761 10912
rect 2825 10848 2841 10912
rect 2905 10848 2921 10912
rect 2985 10848 3001 10912
rect 3065 10848 3073 10912
rect 2753 9824 3073 10848
rect 2753 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2921 9824
rect 2985 9760 3001 9824
rect 3065 9760 3073 9824
rect 2753 8736 3073 9760
rect 4562 12544 4883 13104
rect 4562 12480 4570 12544
rect 4634 12480 4650 12544
rect 4714 12480 4730 12544
rect 4794 12480 4810 12544
rect 4874 12480 4883 12544
rect 4562 11456 4883 12480
rect 4562 11392 4570 11456
rect 4634 11392 4650 11456
rect 4714 11392 4730 11456
rect 4794 11392 4810 11456
rect 4874 11392 4883 11456
rect 4562 10368 4883 11392
rect 4562 10304 4570 10368
rect 4634 10304 4650 10368
rect 4714 10304 4730 10368
rect 4794 10304 4810 10368
rect 4874 10304 4883 10368
rect 4107 9620 4173 9621
rect 4107 9556 4108 9620
rect 4172 9556 4173 9620
rect 4107 9555 4173 9556
rect 2753 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2921 8736
rect 2985 8672 3001 8736
rect 3065 8672 3073 8736
rect 2753 7686 3073 8672
rect 2753 7648 2795 7686
rect 3031 7648 3073 7686
rect 2753 7584 2761 7648
rect 3065 7584 3073 7648
rect 2753 7450 2795 7584
rect 3031 7450 3073 7584
rect 2753 6560 3073 7450
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3073 6560
rect 2753 5472 3073 6496
rect 4110 6493 4170 9555
rect 4562 9499 4883 10304
rect 6372 13088 6692 13104
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 11312 6692 11936
rect 6372 11076 6414 11312
rect 6650 11076 6692 11312
rect 6372 10912 6692 11076
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 5027 9620 5093 9621
rect 5027 9556 5028 9620
rect 5092 9556 5093 9620
rect 5027 9555 5093 9556
rect 4562 9280 4604 9499
rect 4840 9280 4883 9499
rect 4562 9216 4570 9280
rect 4634 9216 4650 9263
rect 4714 9216 4730 9263
rect 4794 9216 4810 9263
rect 4874 9216 4883 9280
rect 4291 8532 4357 8533
rect 4291 8468 4292 8532
rect 4356 8468 4357 8532
rect 4291 8467 4357 8468
rect 4294 7989 4354 8467
rect 4562 8192 4883 9216
rect 4562 8128 4570 8192
rect 4634 8128 4650 8192
rect 4714 8128 4730 8192
rect 4794 8128 4810 8192
rect 4874 8128 4883 8192
rect 4291 7988 4357 7989
rect 4291 7924 4292 7988
rect 4356 7924 4357 7988
rect 4291 7923 4357 7924
rect 4107 6492 4173 6493
rect 4107 6428 4108 6492
rect 4172 6428 4173 6492
rect 4107 6427 4173 6428
rect 4294 5677 4354 7923
rect 4562 7104 4883 8128
rect 4562 7040 4570 7104
rect 4634 7040 4650 7104
rect 4714 7040 4730 7104
rect 4794 7040 4810 7104
rect 4874 7040 4883 7104
rect 4562 6016 4883 7040
rect 5030 6357 5090 9555
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7686 6692 8672
rect 6372 7648 6414 7686
rect 6650 7648 6692 7686
rect 6372 7584 6380 7648
rect 6684 7584 6692 7648
rect 6372 7450 6414 7584
rect 6650 7450 6692 7584
rect 6372 6560 6692 7450
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 5027 6356 5093 6357
rect 5027 6292 5028 6356
rect 5092 6292 5093 6356
rect 5027 6291 5093 6292
rect 4562 5952 4570 6016
rect 4634 5952 4650 6016
rect 4714 5952 4730 6016
rect 4794 5952 4810 6016
rect 4874 5952 4883 6016
rect 4562 5872 4883 5952
rect 4291 5676 4357 5677
rect 4291 5612 4292 5676
rect 4356 5612 4357 5676
rect 4291 5611 4357 5612
rect 4562 5636 4604 5872
rect 4840 5636 4883 5872
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3073 5472
rect 2753 4384 3073 5408
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3073 4384
rect 2753 4059 3073 4320
rect 2753 3823 2795 4059
rect 3031 3823 3073 4059
rect 2753 3296 3073 3823
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3073 3296
rect 2753 2208 3073 3232
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3073 2208
rect 2753 2128 3073 2144
rect 4562 4928 4883 5636
rect 4562 4864 4570 4928
rect 4634 4864 4650 4928
rect 4714 4864 4730 4928
rect 4794 4864 4810 4928
rect 4874 4864 4883 4928
rect 4562 3840 4883 4864
rect 4562 3776 4570 3840
rect 4634 3776 4650 3840
rect 4714 3776 4730 3840
rect 4794 3776 4810 3840
rect 4874 3776 4883 3840
rect 4562 2752 4883 3776
rect 4562 2688 4570 2752
rect 4634 2688 4650 2752
rect 4714 2688 4730 2752
rect 4794 2688 4810 2752
rect 4874 2688 4883 2752
rect 4562 2128 4883 2688
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 4059 6692 4320
rect 6372 3823 6414 4059
rect 6650 3823 6692 4059
rect 6372 3296 6692 3823
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 8181 12544 8501 13104
rect 8181 12480 8189 12544
rect 8253 12480 8269 12544
rect 8333 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8501 12544
rect 8181 11456 8501 12480
rect 8181 11392 8189 11456
rect 8253 11392 8269 11456
rect 8333 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8501 11456
rect 8181 10368 8501 11392
rect 8181 10304 8189 10368
rect 8253 10304 8269 10368
rect 8333 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8501 10368
rect 8181 9499 8501 10304
rect 8181 9280 8223 9499
rect 8459 9280 8501 9499
rect 8181 9216 8189 9280
rect 8253 9216 8269 9263
rect 8333 9216 8349 9263
rect 8413 9216 8429 9263
rect 8493 9216 8501 9280
rect 8181 8192 8501 9216
rect 8181 8128 8189 8192
rect 8253 8128 8269 8192
rect 8333 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8501 8192
rect 8181 7104 8501 8128
rect 8181 7040 8189 7104
rect 8253 7040 8269 7104
rect 8333 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8501 7104
rect 8181 6016 8501 7040
rect 8181 5952 8189 6016
rect 8253 5952 8269 6016
rect 8333 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8501 6016
rect 8181 5872 8501 5952
rect 8181 5636 8223 5872
rect 8459 5636 8501 5872
rect 8181 4928 8501 5636
rect 8181 4864 8189 4928
rect 8253 4864 8269 4928
rect 8333 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8501 4928
rect 8181 3840 8501 4864
rect 8181 3776 8189 3840
rect 8253 3776 8269 3840
rect 8333 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8501 3840
rect 8181 2752 8501 3776
rect 8181 2688 8189 2752
rect 8253 2688 8269 2752
rect 8333 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8501 2752
rect 8181 2128 8501 2688
rect 9990 13088 10311 13104
rect 9990 13024 9998 13088
rect 10062 13024 10078 13088
rect 10142 13024 10158 13088
rect 10222 13024 10238 13088
rect 10302 13024 10311 13088
rect 9990 12000 10311 13024
rect 9990 11936 9998 12000
rect 10062 11936 10078 12000
rect 10142 11936 10158 12000
rect 10222 11936 10238 12000
rect 10302 11936 10311 12000
rect 9990 11312 10311 11936
rect 9990 11076 10032 11312
rect 10268 11076 10311 11312
rect 9990 10912 10311 11076
rect 9990 10848 9998 10912
rect 10062 10848 10078 10912
rect 10142 10848 10158 10912
rect 10222 10848 10238 10912
rect 10302 10848 10311 10912
rect 9990 9824 10311 10848
rect 9990 9760 9998 9824
rect 10062 9760 10078 9824
rect 10142 9760 10158 9824
rect 10222 9760 10238 9824
rect 10302 9760 10311 9824
rect 9990 8736 10311 9760
rect 9990 8672 9998 8736
rect 10062 8672 10078 8736
rect 10142 8672 10158 8736
rect 10222 8672 10238 8736
rect 10302 8672 10311 8736
rect 9990 7686 10311 8672
rect 9990 7648 10032 7686
rect 10268 7648 10311 7686
rect 9990 7584 9998 7648
rect 10302 7584 10311 7648
rect 9990 7450 10032 7584
rect 10268 7450 10311 7584
rect 9990 6560 10311 7450
rect 9990 6496 9998 6560
rect 10062 6496 10078 6560
rect 10142 6496 10158 6560
rect 10222 6496 10238 6560
rect 10302 6496 10311 6560
rect 9990 5472 10311 6496
rect 9990 5408 9998 5472
rect 10062 5408 10078 5472
rect 10142 5408 10158 5472
rect 10222 5408 10238 5472
rect 10302 5408 10311 5472
rect 9990 4384 10311 5408
rect 9990 4320 9998 4384
rect 10062 4320 10078 4384
rect 10142 4320 10158 4384
rect 10222 4320 10238 4384
rect 10302 4320 10311 4384
rect 9990 4059 10311 4320
rect 9990 3823 10032 4059
rect 10268 3823 10311 4059
rect 9990 3296 10311 3823
rect 9990 3232 9998 3296
rect 10062 3232 10078 3296
rect 10142 3232 10158 3296
rect 10222 3232 10238 3296
rect 10302 3232 10311 3296
rect 9990 2208 10311 3232
rect 9990 2144 9998 2208
rect 10062 2144 10078 2208
rect 10142 2144 10158 2208
rect 10222 2144 10238 2208
rect 10302 2144 10311 2208
rect 9990 2128 10311 2144
<< via4 >>
rect 2795 11076 3031 11312
rect 2795 7648 3031 7686
rect 2795 7584 2825 7648
rect 2825 7584 2841 7648
rect 2841 7584 2905 7648
rect 2905 7584 2921 7648
rect 2921 7584 2985 7648
rect 2985 7584 3001 7648
rect 3001 7584 3031 7648
rect 2795 7450 3031 7584
rect 6414 11076 6650 11312
rect 4604 9280 4840 9499
rect 4604 9263 4634 9280
rect 4634 9263 4650 9280
rect 4650 9263 4714 9280
rect 4714 9263 4730 9280
rect 4730 9263 4794 9280
rect 4794 9263 4810 9280
rect 4810 9263 4840 9280
rect 6414 7648 6650 7686
rect 6414 7584 6444 7648
rect 6444 7584 6460 7648
rect 6460 7584 6524 7648
rect 6524 7584 6540 7648
rect 6540 7584 6604 7648
rect 6604 7584 6620 7648
rect 6620 7584 6650 7648
rect 6414 7450 6650 7584
rect 4604 5636 4840 5872
rect 2795 3823 3031 4059
rect 6414 3823 6650 4059
rect 8223 9280 8459 9499
rect 8223 9263 8253 9280
rect 8253 9263 8269 9280
rect 8269 9263 8333 9280
rect 8333 9263 8349 9280
rect 8349 9263 8413 9280
rect 8413 9263 8429 9280
rect 8429 9263 8459 9280
rect 8223 5636 8459 5872
rect 10032 11076 10268 11312
rect 10032 7648 10268 7686
rect 10032 7584 10062 7648
rect 10062 7584 10078 7648
rect 10078 7584 10142 7648
rect 10142 7584 10158 7648
rect 10158 7584 10222 7648
rect 10222 7584 10238 7648
rect 10238 7584 10268 7648
rect 10032 7450 10268 7584
rect 10032 3823 10268 4059
<< metal5 >>
rect 1104 11312 11960 11355
rect 1104 11076 2795 11312
rect 3031 11076 6414 11312
rect 6650 11076 10032 11312
rect 10268 11076 11960 11312
rect 1104 11034 11960 11076
rect 1104 9499 11960 9541
rect 1104 9263 4604 9499
rect 4840 9263 8223 9499
rect 8459 9263 11960 9499
rect 1104 9221 11960 9263
rect 1104 7686 11960 7728
rect 1104 7450 2795 7686
rect 3031 7450 6414 7686
rect 6650 7450 10032 7686
rect 10268 7450 11960 7686
rect 1104 7408 11960 7450
rect 1104 5872 11960 5915
rect 1104 5636 4604 5872
rect 4840 5636 8223 5872
rect 8459 5636 11960 5872
rect 1104 5594 11960 5636
rect 1104 4059 11960 4101
rect 1104 3823 2795 4059
rect 3031 3823 6414 4059
rect 6650 3823 10032 4059
rect 10268 3823 11960 4059
rect 1104 3781 11960 3823
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1619947793
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12
timestamp 1619947793
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1619947793
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1619947793
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _159_
timestamp 1619947793
transform 1 0 1932 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _141_
timestamp 1619947793
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1619947793
transform 1 0 4784 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1619947793
transform 1 0 3680 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39
timestamp 1619947793
transform 1 0 4692 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1619947793
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24
timestamp 1619947793
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1619947793
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _146_
timestamp 1619947793
transform 1 0 4048 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1619947793
transform 1 0 6808 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1619947793
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1619947793
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1619947793
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1619947793
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _132_
timestamp 1619947793
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _111_
timestamp 1619947793
transform 1 0 5428 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1619947793
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1619947793
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _161_
timestamp 1619947793
transform 1 0 7728 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _103_
timestamp 1619947793
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1619947793
transform 1 0 10212 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1619947793
transform 1 0 9476 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1619947793
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1619947793
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _112_
timestamp 1619947793
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _097_
timestamp 1619947793
transform 1 0 10304 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_107
timestamp 1619947793
transform 1 0 10948 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114
timestamp 1619947793
transform 1 0 11592 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106
timestamp 1619947793
transform 1 0 10856 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1619947793
transform -1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1619947793
transform -1 0 11960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_12
timestamp 1619947793
transform 1 0 2208 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1619947793
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1619947793
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1619947793
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _093_
timestamp 1619947793
transform 1 0 1564 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1619947793
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1619947793
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1619947793
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1619947793
transform 1 0 5980 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1619947793
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _078_
timestamp 1619947793
transform 1 0 5336 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _155_
timestamp 1619947793
transform 1 0 7084 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_2_102
timestamp 1619947793
transform 1 0 10488 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1619947793
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1619947793
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _084_
timestamp 1619947793
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_114
timestamp 1619947793
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1619947793
transform -1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_16
timestamp 1619947793
transform 1 0 2576 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1619947793
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1619947793
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _115_
timestamp 1619947793
transform 1 0 1932 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1619947793
transform 1 0 4784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_28
timestamp 1619947793
transform 1 0 3680 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1619947793
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1619947793
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _162_
timestamp 1619947793
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _098_
timestamp 1619947793
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1619947793
transform 1 0 8556 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1619947793
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _136_
timestamp 1619947793
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_114
timestamp 1619947793
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1619947793
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1619947793
transform -1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 1619947793
transform 1 0 2576 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1619947793
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _142_
timestamp 1619947793
transform 1 0 1380 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_4_39
timestamp 1619947793
transform 1 0 4692 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1619947793
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1619947793
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _081_
timestamp 1619947793
transform 1 0 4048 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp 1619947793
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _153_
timestamp 1619947793
transform 1 0 5704 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1619947793
transform 1 0 7452 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _102_
timestamp 1619947793
transform 1 0 8188 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_4_102
timestamp 1619947793
transform 1 0 10488 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_84
timestamp 1619947793
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1619947793
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _117_
timestamp 1619947793
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_114
timestamp 1619947793
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1619947793
transform -1 0 11960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1619947793
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_12
timestamp 1619947793
transform 1 0 2208 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1619947793
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _083_
timestamp 1619947793
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1619947793
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_24
timestamp 1619947793
transform 1 0 3312 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1619947793
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _114_
timestamp 1619947793
transform 1 0 4048 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1619947793
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1619947793
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1619947793
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1619947793
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1619947793
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_66
timestamp 1619947793
transform 1 0 7176 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _157_
timestamp 1619947793
transform 1 0 7912 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1619947793
transform 1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1619947793
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1619947793
transform 1 0 9660 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1619947793
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_107
timestamp 1619947793
transform 1 0 10948 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1619947793
transform -1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1619947793
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1619947793
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_19
timestamp 1619947793
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1619947793
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1619947793
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1619947793
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1619947793
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1619947793
transform 1 0 1472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_36
timestamp 1619947793
transform 1 0 4416 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1619947793
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _145_
timestamp 1619947793
transform 1 0 4048 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _128_
timestamp 1619947793
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1619947793
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_46
timestamp 1619947793
transform 1 0 5336 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_44
timestamp 1619947793
transform 1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_50
timestamp 1619947793
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _119_
timestamp 1619947793
transform 1 0 6440 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1619947793
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1619947793
transform 1 0 6072 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1619947793
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1619947793
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1619947793
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_75
timestamp 1619947793
transform 1 0 8004 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_67
timestamp 1619947793
transform 1 0 7268 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _120_
timestamp 1619947793
transform 1 0 7360 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _082_
timestamp 1619947793
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_99
timestamp 1619947793
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_102
timestamp 1619947793
transform 1 0 10488 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1619947793
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1619947793
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _100_
timestamp 1619947793
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _087_
timestamp 1619947793
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_111
timestamp 1619947793
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_114
timestamp 1619947793
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1619947793
transform -1 0 11960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1619947793
transform -1 0 11960 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1619947793
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1619947793
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1619947793
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1619947793
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1619947793
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1619947793
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1619947793
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1619947793
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_4  _140_
timestamp 1619947793
transform 1 0 4784 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_58
timestamp 1619947793
transform 1 0 6440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_69
timestamp 1619947793
transform 1 0 7452 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1619947793
transform 1 0 7176 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _095_
timestamp 1619947793
transform 1 0 8188 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1619947793
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1619947793
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1619947793
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _116_
timestamp 1619947793
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1619947793
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1619947793
transform -1 0 11960 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1619947793
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_12
timestamp 1619947793
transform 1 0 2208 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1619947793
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1619947793
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1619947793
transform 1 0 1932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_29
timestamp 1619947793
transform 1 0 3772 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1619947793
transform 1 0 4876 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_4  _123_
timestamp 1619947793
transform 1 0 3128 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_9_62
timestamp 1619947793
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1619947793
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_82
timestamp 1619947793
transform 1 0 8648 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_68
timestamp 1619947793
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _106_
timestamp 1619947793
transform 1 0 7452 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1619947793
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _134_
timestamp 1619947793
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1619947793
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1619947793
transform -1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1619947793
transform 1 0 2300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1619947793
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1619947793
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _131_
timestamp 1619947793
transform 1 0 1472 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1619947793
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1619947793
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _124_
timestamp 1619947793
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _107_
timestamp 1619947793
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1619947793
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _158_
timestamp 1619947793
transform 1 0 5888 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1619947793
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_71
timestamp 1619947793
transform 1 0 7636 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1619947793
transform 1 0 8372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_102
timestamp 1619947793
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1619947793
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1619947793
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _137_
timestamp 1619947793
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1619947793
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1619947793
transform -1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_19
timestamp 1619947793
transform 1 0 2852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1619947793
transform 1 0 1748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1619947793
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1619947793
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_41
timestamp 1619947793
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_33
timestamp 1619947793
transform 1 0 4140 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1619947793
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1619947793
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1619947793
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1619947793
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1619947793
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _143_
timestamp 1619947793
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1619947793
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1619947793
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1619947793
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1619947793
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _160_
timestamp 1619947793
transform 1 0 9200 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_11_107
timestamp 1619947793
transform 1 0 10948 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1619947793
transform -1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1619947793
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _151_
timestamp 1619947793
transform 1 0 1380 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_38
timestamp 1619947793
transform 1 0 4600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1619947793
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1619947793
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1619947793
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1619947793
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1619947793
transform 1 0 4232 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_62
timestamp 1619947793
transform 1 0 6808 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_50
timestamp 1619947793
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_76
timestamp 1619947793
transform 1 0 8096 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_70
timestamp 1619947793
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1619947793
transform 1 0 7820 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1619947793
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1619947793
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1619947793
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1619947793
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _089_
timestamp 1619947793
transform 1 0 10304 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_107
timestamp 1619947793
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1619947793
transform -1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1619947793
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1619947793
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1619947793
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1619947793
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1619947793
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1619947793
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1619947793
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _139_
timestamp 1619947793
transform 1 0 1840 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _126_
timestamp 1619947793
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1619947793
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1619947793
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1619947793
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _149_
timestamp 1619947793
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _122_
timestamp 1619947793
transform 1 0 4048 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_14_61
timestamp 1619947793
transform 1 0 6716 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_46
timestamp 1619947793
transform 1 0 5336 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1619947793
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1619947793
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1619947793
transform 1 0 5520 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1619947793
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1619947793
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _148_
timestamp 1619947793
transform 1 0 6072 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1619947793
transform 1 0 8464 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_72
timestamp 1619947793
transform 1 0 7728 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1619947793
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_74
timestamp 1619947793
transform 1 0 7912 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1619947793
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1619947793
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _121_
timestamp 1619947793
transform 1 0 8740 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1619947793
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1619947793
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1619947793
transform 1 0 10580 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_95
timestamp 1619947793
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1619947793
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _109_
timestamp 1619947793
transform 1 0 9844 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1619947793
transform 1 0 10672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_107
timestamp 1619947793
transform 1 0 10948 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_107
timestamp 1619947793
transform 1 0 10948 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1619947793
transform -1 0 11960 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1619947793
transform -1 0 11960 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1619947793
transform 1 0 2484 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1619947793
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1619947793
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1619947793
transform 1 0 4784 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _150_
timestamp 1619947793
transform 1 0 3036 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1619947793
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_52
timestamp 1619947793
transform 1 0 5888 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1619947793
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1619947793
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_77
timestamp 1619947793
transform 1 0 8188 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_65
timestamp 1619947793
transform 1 0 7084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _154_
timestamp 1619947793
transform 1 0 8740 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_102
timestamp 1619947793
transform 1 0 10488 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_114
timestamp 1619947793
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1619947793
transform -1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1619947793
transform 1 0 2392 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1619947793
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1619947793
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _130_
timestamp 1619947793
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1619947793
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1619947793
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1619947793
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _152_
timestamp 1619947793
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1619947793
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _156_
timestamp 1619947793
transform 1 0 6532 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_78
timestamp 1619947793
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1619947793
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1619947793
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1619947793
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _138_
timestamp 1619947793
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1619947793
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1619947793
transform -1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1619947793
transform 1 0 2484 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1619947793
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1619947793
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1619947793
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_23
timestamp 1619947793
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _099_
timestamp 1619947793
transform 1 0 3312 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1619947793
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1619947793
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1619947793
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _118_
timestamp 1619947793
transform 1 0 5336 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_79
timestamp 1619947793
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _133_
timestamp 1619947793
transform 1 0 7544 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_102
timestamp 1619947793
transform 1 0 10488 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1619947793
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _085_
timestamp 1619947793
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_114
timestamp 1619947793
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1619947793
transform -1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_19
timestamp 1619947793
transform 1 0 2852 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1619947793
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1619947793
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1619947793
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _147_
timestamp 1619947793
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1619947793
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1619947793
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1619947793
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _105_
timestamp 1619947793
transform 1 0 4876 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1619947793
transform 1 0 5980 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1619947793
transform 1 0 7084 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _101_
timestamp 1619947793
transform 1 0 7636 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1619947793
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1619947793
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1619947793
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1619947793
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_105
timestamp 1619947793
transform 1 0 10764 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1619947793
transform -1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1619947793
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1619947793
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1619947793
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_41
timestamp 1619947793
transform 1 0 4876 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1619947793
transform 1 0 3588 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1619947793
transform 1 0 3956 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _113_
timestamp 1619947793
transform 1 0 4048 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1619947793
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1619947793
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1619947793
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_75
timestamp 1619947793
transform 1 0 8004 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_63
timestamp 1619947793
transform 1 0 6900 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1619947793
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 1619947793
transform 1 0 9108 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1619947793
transform 1 0 9660 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_114
timestamp 1619947793
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1619947793
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1619947793
transform -1 0 11960 0 1 12512
box -38 -48 314 592
<< labels >>
rlabel metal3 s 12902 10616 13102 10736 4 change[0]
port 1 nsew
rlabel metal3 s 12902 13608 13102 13728 4 change[1]
port 2 nsew
rlabel metal3 s 0 1504 200 1624 4 choice[0]
port 3 nsew
rlabel metal3 s 0 4496 200 4616 4 choice[1]
port 4 nsew
rlabel metal3 s 0 7488 200 7608 4 choice[2]
port 5 nsew
rlabel metal2 s 3238 0 3294 200 4 clk
port 6 nsew
rlabel metal3 s 0 10616 200 10736 4 coin[0]
port 7 nsew
rlabel metal3 s 0 13608 200 13728 4 coin[1]
port 8 nsew
rlabel metal3 s 12902 1504 13102 1624 4 out[0]
port 9 nsew
rlabel metal3 s 12902 4496 13102 4616 4 out[1]
port 10 nsew
rlabel metal3 s 12902 7488 13102 7608 4 out[2]
port 11 nsew
rlabel metal2 s 9770 0 9826 200 4 reset
port 12 nsew
rlabel metal4 s 9991 2128 10311 13104 4 VPWR
port 13 nsew
rlabel metal4 s 6372 2128 6692 13104 4 VPWR
port 13 nsew
rlabel metal4 s 2753 2128 3073 13104 4 VPWR
port 13 nsew
rlabel metal5 s 1104 11035 11960 11355 4 VPWR
port 13 nsew
rlabel metal5 s 1104 7408 11960 7728 4 VPWR
port 13 nsew
rlabel metal5 s 1104 3781 11960 4101 4 VPWR
port 13 nsew
rlabel metal4 s 8181 2128 8501 13104 4 VGND
port 14 nsew
rlabel metal4 s 4563 2128 4883 13104 4 VGND
port 14 nsew
rlabel metal5 s 1104 9221 11960 9541 4 VGND
port 14 nsew
rlabel metal5 s 1104 5595 11960 5915 4 VGND
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 13102 13728
<< end >>
