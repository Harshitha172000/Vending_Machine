* NGSPICE file created from vm.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt vm change[0] change[1] choice[0] choice[1] choice[2] clk coin[0] coin[1] out[0]
+ out[1] out[2] reset VPWR VGND
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_131_ _129_/Y choice[1] _130_/X _125_/Y VGND VGND VPWR VPWR _131_/X sky130_fd_sc_hd__and4_4
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_114_ _079_/Y _114_/B VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__and2_4
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_130_ _130_/A _085_/C _126_/X VGND VGND VPWR VPWR _130_/X sky130_fd_sc_hd__and3_4
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_113_ _113_/A _113_/B _113_/C VGND VGND VPWR VPWR _114_/B sky130_fd_sc_hd__or3_4
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_112_ _137_/D _111_/X _147_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__o21a_4
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ _113_/B _133_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__and2_4
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_110_ _152_/Q VGND VGND VPWR VPWR _113_/B sky130_fd_sc_hd__buf_2
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _147_/C _138_/D _098_/X _148_/A VGND VGND VPWR VPWR _100_/C sky130_fd_sc_hd__a211o_4
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_098_ _147_/A _147_/B _098_/C VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__and3_4
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_097_ _080_/X _081_/X VGND VGND VPWR VPWR _098_/C sky130_fd_sc_hd__or2_4
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_149_ _149_/A _146_/X _149_/C VGND VGND VPWR VPWR _162_/D sky130_fd_sc_hd__and3_4
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ _148_/A _148_/B VGND VGND VPWR VPWR _149_/C sky130_fd_sc_hd__or2_4
X_096_ _143_/B VGND VGND VPWR VPWR _147_/A sky130_fd_sc_hd__inv_2
X_079_ _078_/X VGND VGND VPWR VPWR _079_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ coin[0] _092_/A VGND VGND VPWR VPWR _143_/B sky130_fd_sc_hd__and2_4
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_147_ _147_/A _147_/B _147_/C VGND VGND VPWR VPWR _148_/B sky130_fd_sc_hd__and3_4
X_078_ coin[0] coin[1] VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__or2_4
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_094_ _147_/B VGND VGND VPWR VPWR _138_/D sky130_fd_sc_hd__inv_2
X_129_ choice[2] VGND VGND VPWR VPWR _129_/Y sky130_fd_sc_hd__inv_2
X_077_ _133_/C VGND VGND VPWR VPWR _149_/A sky130_fd_sc_hd__buf_2
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_146_ change[1] _088_/Y VGND VGND VPWR VPWR _146_/X sky130_fd_sc_hd__or2_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_093_ _133_/A _133_/B VGND VGND VPWR VPWR _147_/B sky130_fd_sc_hd__or2_4
X_162_ _157_/CLK _162_/D VGND VGND VPWR VPWR change[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_076_ _130_/A VGND VGND VPWR VPWR _133_/C sky130_fd_sc_hd__buf_2
X_145_ _130_/X _140_/X _141_/X _144_/Y VGND VGND VPWR VPWR _145_/X sky130_fd_sc_hd__a211o_4
X_128_ _149_/A _085_/C _127_/Y VGND VGND VPWR VPWR _128_/X sky130_fd_sc_hd__and3_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ _092_/A VGND VGND VPWR VPWR _133_/B sky130_fd_sc_hd__buf_2
X_161_ _157_/CLK _161_/D VGND VGND VPWR VPWR change[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_144_ _143_/X VGND VGND VPWR VPWR _144_/Y sky130_fd_sc_hd__inv_2
X_075_ reset VGND VGND VPWR VPWR _130_/A sky130_fd_sc_hd__inv_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_127_ _126_/X VGND VGND VPWR VPWR _127_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_160_ _154_/CLK _160_/D VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__dfxtp_4
X_143_ reset _143_/B _142_/Y VGND VGND VPWR VPWR _143_/X sky130_fd_sc_hd__or3_4
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ coin[1] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__inv_2
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_126_ choice[2] choice[1] _125_/Y VGND VGND VPWR VPWR _126_/X sky130_fd_sc_hd__or3_4
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _085_/X _078_/X out[1] VGND VGND VPWR VPWR _117_/B sky130_fd_sc_hd__a21o_4
X_090_ coin[0] VGND VGND VPWR VPWR _133_/A sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_125_ choice[0] VGND VGND VPWR VPWR _125_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_142_ _113_/B _147_/B _081_/X VGND VGND VPWR VPWR _142_/Y sky130_fd_sc_hd__a21oi_4
X_108_ _107_/X VGND VGND VPWR VPWR _160_/D sky130_fd_sc_hd__inv_2
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_141_ _113_/A _116_/A reset _102_/X VGND VGND VPWR VPWR _141_/X sky130_fd_sc_hd__or4_4
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ _149_/A _124_/B _123_/X VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__and3_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_107_ reset _107_/B _107_/C VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__or3_4
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_140_ _129_/Y choice[1] choice[0] choice[2] _135_/Y VGND VGND VPWR VPWR _140_/X sky130_fd_sc_hd__o32a_4
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_106_ _080_/X _118_/B out[2] VGND VGND VPWR VPWR _107_/C sky130_fd_sc_hd__a21oi_4
X_123_ _123_/A _123_/B VGND VGND VPWR VPWR _123_/X sky130_fd_sc_hd__or2_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _154_/CLK sky130_fd_sc_hd__clkbuf_1
X_122_ _113_/A _121_/X out[0] _078_/X VGND VGND VPWR VPWR _123_/B sky130_fd_sc_hd__o22a_4
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_105_ _143_/B _101_/Y _118_/B VGND VGND VPWR VPWR _107_/B sky130_fd_sc_hd__o21a_4
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_121_ _113_/C _120_/X _147_/A VGND VGND VPWR VPWR _121_/X sky130_fd_sc_hd__o21a_4
X_104_ _104_/A VGND VGND VPWR VPWR _118_/B sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _157_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_120_ _092_/A _119_/X VGND VGND VPWR VPWR _120_/X sky130_fd_sc_hd__and2_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_103_ _102_/X _079_/Y _086_/Y VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__a21o_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_102_ _085_/A _080_/X VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__or2_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ _133_/B _084_/X _080_/X VGND VGND VPWR VPWR _101_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_100_ _149_/A _100_/B _100_/C VGND VGND VPWR VPWR _161_/D sky130_fd_sc_hd__and3_4
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_159_ _157_/CLK _159_/D VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ change[0] _088_/Y VGND VGND VPWR VPWR _100_/B sky130_fd_sc_hd__or2_4
X_158_ _154_/CLK _124_/X VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ _148_/A VGND VGND VPWR VPWR _088_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_157_ _157_/CLK _136_/X VGND VGND VPWR VPWR _085_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_156_ _154_/CLK _134_/X VGND VGND VPWR VPWR _085_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_087_ _079_/Y _083_/X _086_/Y VGND VGND VPWR VPWR _148_/A sky130_fd_sc_hd__a21o_4
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_139_ _137_/X _139_/B VGND VGND VPWR VPWR _153_/D sky130_fd_sc_hd__or2_4
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_155_ _157_/CLK _132_/X VGND VGND VPWR VPWR _137_/D sky130_fd_sc_hd__dfxtp_4
X_086_ _085_/X VGND VGND VPWR VPWR _086_/Y sky130_fd_sc_hd__inv_2
X_138_ _133_/C _147_/A _113_/B _138_/D VGND VGND VPWR VPWR _139_/B sky130_fd_sc_hd__and4_4
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ _085_/A _085_/B _085_/C _084_/X VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__or4_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_154_ _154_/CLK _128_/X VGND VGND VPWR VPWR _113_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_137_ _133_/A _133_/B _133_/C _137_/D VGND VGND VPWR VPWR _137_/X sky130_fd_sc_hd__and4_4
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_084_ _113_/A _116_/A _152_/Q _081_/X VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__or4_4
X_136_ choice[2] _135_/Y _125_/Y _130_/X VGND VGND VPWR VPWR _136_/X sky130_fd_sc_hd__and4_4
X_153_ _157_/CLK _153_/D VGND VGND VPWR VPWR _116_/A sky130_fd_sc_hd__dfxtp_4
X_119_ _152_/Q _116_/A _137_/D VGND VGND VPWR VPWR _119_/X sky130_fd_sc_hd__or3_4
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ _154_/CLK _131_/X VGND VGND VPWR VPWR _152_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ _080_/X _081_/X _152_/Q _147_/C VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__or4_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_118_ out[0] _118_/B VGND VGND VPWR VPWR _124_/B sky130_fd_sc_hd__or2_4
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_135_ choice[1] VGND VGND VPWR VPWR _135_/Y sky130_fd_sc_hd__inv_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_151_ _154_/CLK _151_/D VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__dfxtp_4
X_134_ _129_/Y choice[1] _130_/X choice[0] VGND VGND VPWR VPWR _134_/X sky130_fd_sc_hd__and4_4
X_082_ _113_/A _116_/A _085_/A VGND VGND VPWR VPWR _147_/C sky130_fd_sc_hd__or3_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_117_ _149_/A _117_/B _117_/C VGND VGND VPWR VPWR _159_/D sky130_fd_sc_hd__and3_4
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_150_ _154_/CLK _145_/X VGND VGND VPWR VPWR _085_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ _113_/C _137_/D VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__or2_4
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_133_ _133_/A _133_/B _133_/C _113_/C VGND VGND VPWR VPWR _151_/D sky130_fd_sc_hd__and4_4
XFILLER_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ _116_/A _112_/X _114_/X _123_/A VGND VGND VPWR VPWR _117_/C sky130_fd_sc_hd__or4_4
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_080_ _085_/B VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__buf_2
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_132_ _133_/A _133_/B _133_/C _113_/B VGND VGND VPWR VPWR _132_/X sky130_fd_sc_hd__and4_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_115_ _085_/A _104_/A VGND VGND VPWR VPWR _123_/A sky130_fd_sc_hd__or2_4
.ends

