module vm (clk,
    reset,
    VPWR,
    VGND,
    change,
    choice,
    coin,
    out);
 input clk;
 input reset;
 input VPWR;
 input VGND;
 output [1:0] change;
 input [2:0] choice;
 input [1:0] coin;
 output [2:0] out;

 sky130_fd_sc_hd__inv_2 _075_ (.A(reset),
    .Y(_019_));
 sky130_fd_sc_hd__buf_2 _076_ (.A(_019_),
    .X(_020_));
 sky130_fd_sc_hd__buf_2 _077_ (.A(_020_),
    .X(_021_));
 sky130_fd_sc_hd__or2_4 _078_ (.A(coin[0]),
    .B(coin[1]),
    .X(_022_));
 sky130_fd_sc_hd__inv_2 _079_ (.A(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__buf_2 _080_ (.A(\state[7] ),
    .X(_024_));
 sky130_fd_sc_hd__or2_4 _081_ (.A(\state[4] ),
    .B(\state[5] ),
    .X(_025_));
 sky130_fd_sc_hd__or3_4 _082_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(\state[6] ),
    .X(_026_));
 sky130_fd_sc_hd__or4_4 _083_ (.A(_024_),
    .B(_025_),
    .C(\state[2] ),
    .D(_026_),
    .X(_027_));
 sky130_fd_sc_hd__or4_4 _084_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(\state[2] ),
    .D(_025_),
    .X(_028_));
 sky130_fd_sc_hd__or4_4 _085_ (.A(\state[6] ),
    .B(\state[7] ),
    .C(\state[0] ),
    .D(_028_),
    .X(_029_));
 sky130_fd_sc_hd__inv_2 _086_ (.A(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__a21o_4 _087_ (.A1(_023_),
    .A2(_027_),
    .B1(_030_),
    .X(_031_));
 sky130_fd_sc_hd__inv_2 _088_ (.A(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__or2_4 _089_ (.A(change[0]),
    .B(_032_),
    .X(_033_));
 sky130_fd_sc_hd__buf_2 _090_ (.A(coin[0]),
    .X(_034_));
 sky130_fd_sc_hd__inv_2 _091_ (.A(coin[1]),
    .Y(_035_));
 sky130_fd_sc_hd__buf_2 _092_ (.A(_035_),
    .X(_036_));
 sky130_fd_sc_hd__or2_4 _093_ (.A(_034_),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__inv_2 _094_ (.A(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__and2_4 _095_ (.A(coin[0]),
    .B(_035_),
    .X(_039_));
 sky130_fd_sc_hd__inv_2 _096_ (.A(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__or2_4 _097_ (.A(_024_),
    .B(_025_),
    .X(_041_));
 sky130_fd_sc_hd__and3_4 _098_ (.A(_040_),
    .B(_037_),
    .C(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a211o_4 _099_ (.A1(_026_),
    .A2(_038_),
    .B1(_042_),
    .C1(_031_),
    .X(_043_));
 sky130_fd_sc_hd__and3_4 _100_ (.A(_021_),
    .B(_033_),
    .C(_043_),
    .X(_011_));
 sky130_fd_sc_hd__a21oi_4 _101_ (.A1(_036_),
    .A2(_028_),
    .B1(_024_),
    .Y(_044_));
 sky130_fd_sc_hd__or2_4 _102_ (.A(\state[6] ),
    .B(_024_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_4 _103_ (.A1(_045_),
    .A2(_023_),
    .B1(_030_),
    .X(_046_));
 sky130_fd_sc_hd__inv_2 _104_ (.A(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__o21a_4 _105_ (.A1(_039_),
    .A2(_044_),
    .B1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__a21oi_4 _106_ (.A1(_024_),
    .A2(_047_),
    .B1(out[2]),
    .Y(_049_));
 sky130_fd_sc_hd__or3_4 _107_ (.A(reset),
    .B(_048_),
    .C(_049_),
    .X(_050_));
 sky130_fd_sc_hd__inv_2 _108_ (.A(_050_),
    .Y(_010_));
 sky130_fd_sc_hd__a21o_4 _109_ (.A1(_029_),
    .A2(_022_),
    .B1(out[1]),
    .X(_051_));
 sky130_fd_sc_hd__buf_2 _110_ (.A(\state[2] ),
    .X(_052_));
 sky130_fd_sc_hd__and2_4 _111_ (.A(_052_),
    .B(_034_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_4 _112_ (.A1(\state[5] ),
    .A2(_053_),
    .B1(_040_),
    .X(_054_));
 sky130_fd_sc_hd__or3_4 _113_ (.A(\state[1] ),
    .B(_052_),
    .C(\state[4] ),
    .X(_055_));
 sky130_fd_sc_hd__and2_4 _114_ (.A(_023_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__or2_4 _115_ (.A(\state[6] ),
    .B(_046_),
    .X(_057_));
 sky130_fd_sc_hd__or4_4 _116_ (.A(\state[3] ),
    .B(_054_),
    .C(_056_),
    .D(_057_),
    .X(_058_));
 sky130_fd_sc_hd__and3_4 _117_ (.A(_021_),
    .B(_051_),
    .C(_058_),
    .X(_009_));
 sky130_fd_sc_hd__or2_4 _118_ (.A(out[0]),
    .B(_047_),
    .X(_059_));
 sky130_fd_sc_hd__or3_4 _119_ (.A(\state[2] ),
    .B(\state[3] ),
    .C(\state[5] ),
    .X(_060_));
 sky130_fd_sc_hd__and2_4 _120_ (.A(_035_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__o21a_4 _121_ (.A1(\state[4] ),
    .A2(_061_),
    .B1(_040_),
    .X(_062_));
 sky130_fd_sc_hd__o22a_4 _122_ (.A1(\state[1] ),
    .A2(_062_),
    .B1(out[0]),
    .B2(_022_),
    .X(_063_));
 sky130_fd_sc_hd__or2_4 _123_ (.A(_057_),
    .B(_063_),
    .X(_064_));
 sky130_fd_sc_hd__and3_4 _124_ (.A(_021_),
    .B(_059_),
    .C(_064_),
    .X(_008_));
 sky130_fd_sc_hd__inv_2 _125_ (.A(choice[0]),
    .Y(_065_));
 sky130_fd_sc_hd__or3_4 _126_ (.A(choice[2]),
    .B(choice[1]),
    .C(_065_),
    .X(_066_));
 sky130_fd_sc_hd__inv_2 _127_ (.A(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__and3_4 _128_ (.A(_021_),
    .B(\state[0] ),
    .C(_067_),
    .X(_002_));
 sky130_fd_sc_hd__inv_2 _129_ (.A(choice[2]),
    .Y(_068_));
 sky130_fd_sc_hd__and3_4 _130_ (.A(_019_),
    .B(\state[0] ),
    .C(_066_),
    .X(_069_));
 sky130_fd_sc_hd__and4_4 _131_ (.A(_068_),
    .B(choice[1]),
    .C(_069_),
    .D(_065_),
    .X(_001_));
 sky130_fd_sc_hd__and4_4 _132_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(_052_),
    .X(_003_));
 sky130_fd_sc_hd__and4_4 _133_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(\state[4] ),
    .X(_000_));
 sky130_fd_sc_hd__and4_4 _134_ (.A(_068_),
    .B(choice[1]),
    .C(_069_),
    .D(choice[0]),
    .X(_004_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(choice[1]),
    .Y(_070_));
 sky130_fd_sc_hd__and4_4 _136_ (.A(choice[2]),
    .B(_070_),
    .C(_065_),
    .D(_069_),
    .X(_005_));
 sky130_fd_sc_hd__and4_4 _137_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(\state[5] ),
    .X(_071_));
 sky130_fd_sc_hd__and4_4 _138_ (.A(_020_),
    .B(_040_),
    .C(_052_),
    .D(_038_),
    .X(_072_));
 sky130_fd_sc_hd__or2_4 _139_ (.A(_071_),
    .B(_072_),
    .X(_007_));
 sky130_fd_sc_hd__o32a_4 _140_ (.A1(_068_),
    .A2(choice[1]),
    .A3(choice[0]),
    .B1(choice[2]),
    .B2(_070_),
    .X(_073_));
 sky130_fd_sc_hd__or4_4 _141_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(reset),
    .D(_045_),
    .X(_074_));
 sky130_fd_sc_hd__a21oi_4 _142_ (.A1(_052_),
    .A2(_037_),
    .B1(_025_),
    .Y(_013_));
 sky130_fd_sc_hd__or3_4 _143_ (.A(reset),
    .B(_039_),
    .C(_013_),
    .X(_014_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__a211o_4 _145_ (.A1(_069_),
    .A2(_073_),
    .B1(_074_),
    .C1(_015_),
    .X(_006_));
 sky130_fd_sc_hd__or2_4 _146_ (.A(change[1]),
    .B(_032_),
    .X(_016_));
 sky130_fd_sc_hd__and3_4 _147_ (.A(_040_),
    .B(_037_),
    .C(_026_),
    .X(_017_));
 sky130_fd_sc_hd__or2_4 _148_ (.A(_031_),
    .B(_017_),
    .X(_018_));
 sky130_fd_sc_hd__and3_4 _149_ (.A(_021_),
    .B(_016_),
    .C(_018_),
    .X(_012_));
 sky130_fd_sc_hd__dfxtp_4 _150_ (.D(_006_),
    .Q(\state[0] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _151_ (.D(_000_),
    .Q(\state[1] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _152_ (.D(_001_),
    .Q(\state[2] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _153_ (.D(_007_),
    .Q(\state[3] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _154_ (.D(_002_),
    .Q(\state[4] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _155_ (.D(_003_),
    .Q(\state[5] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _156_ (.D(_004_),
    .Q(\state[6] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _157_ (.D(_005_),
    .Q(\state[7] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _158_ (.D(_008_),
    .Q(out[0]),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _159_ (.D(_009_),
    .Q(out[1]),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _160_ (.D(_010_),
    .Q(out[2]),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _161_ (.D(_011_),
    .Q(change[0]),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _162_ (.D(_012_),
    .Q(change[1]),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_210 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_107 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_133 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_160 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_49 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_19 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_126 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_19 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_39 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_170 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_95 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_112 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_82 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_210 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_112 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_160 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_101 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_60 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_43 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_67 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_22 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_34 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_60 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_216 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_71 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_95 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_210 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_179 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_12 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_36 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_210 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_95 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_217 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_214 ();
endmodule
