VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vm
  CLASS BLOCK ;
  FOREIGN vm ;
  ORIGIN 0.000 0.000 ;
  SIZE 65.510 BY 68.640 ;
  PIN change[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.510 53.080 65.510 53.680 ;
    END
  END change[0]
  PIN change[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.510 68.040 65.510 68.640 ;
    END
  END change[1]
  PIN choice[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 1.000 8.120 ;
    END
  END choice[0]
  PIN choice[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 1.000 23.080 ;
    END
  END choice[1]
  PIN choice[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 1.000 38.040 ;
    END
  END choice[2]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 1.000 ;
    END
  END clk
  PIN coin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 1.000 53.680 ;
    END
  END coin[0]
  PIN coin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 1.000 68.640 ;
    END
  END coin[1]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.510 7.520 65.510 8.120 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.510 22.480 65.510 23.080 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.510 37.440 65.510 38.040 ;
    END
  END out[2]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 1.000 ;
    END
  END reset
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 49.955 10.640 51.555 65.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.860 10.640 33.460 65.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.765 10.640 15.365 65.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 55.175 59.800 56.775 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 37.040 59.800 38.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 18.905 59.800 20.505 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 40.905 10.640 42.505 65.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 22.815 10.640 24.415 65.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 46.105 59.800 47.705 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 27.975 59.800 29.575 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 59.800 65.365 ;
      LAYER met1 ;
        RECT 5.520 9.560 59.800 65.520 ;
      LAYER met2 ;
        RECT 6.990 1.280 55.110 68.525 ;
        RECT 6.990 1.000 15.910 1.280 ;
        RECT 16.750 1.000 48.570 1.280 ;
        RECT 49.410 1.000 55.110 1.280 ;
      LAYER met3 ;
        RECT 1.400 67.640 64.110 68.505 ;
        RECT 1.000 54.080 64.510 67.640 ;
        RECT 1.400 52.680 64.110 54.080 ;
        RECT 1.000 38.440 64.510 52.680 ;
        RECT 1.400 37.040 64.110 38.440 ;
        RECT 1.000 23.480 64.510 37.040 ;
        RECT 1.400 22.080 64.110 23.480 ;
        RECT 1.000 8.520 64.510 22.080 ;
        RECT 1.400 7.655 64.110 8.520 ;
      LAYER met4 ;
        RECT 20.535 10.640 22.415 65.520 ;
        RECT 24.815 10.640 31.460 65.520 ;
        RECT 33.860 10.640 40.505 65.520 ;
        RECT 42.905 10.640 49.555 65.520 ;
      LAYER met5 ;
        RECT 5.520 49.305 59.800 53.575 ;
        RECT 5.520 40.240 59.800 44.505 ;
        RECT 5.520 31.175 59.800 35.440 ;
  END
END vm
END LIBRARY

