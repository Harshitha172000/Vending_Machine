magic
tech sky130A
magscale 1 2
timestamp 1617727117
<< obsli1 >>
rect 1104 2159 21436 22321
<< obsm1 >>
rect 566 2128 21974 22352
<< metal2 >>
rect 3330 23933 3386 24733
rect 9586 23933 9642 24733
rect 15842 23933 15898 24733
rect 21914 23933 21970 24733
rect 570 0 626 800
rect 6642 0 6698 800
rect 12898 0 12954 800
rect 19154 0 19210 800
<< obsm2 >>
rect 572 23877 3274 23933
rect 3442 23877 9530 23933
rect 9698 23877 15786 23933
rect 15954 23877 21858 23933
rect 572 856 21968 23877
rect 682 800 6586 856
rect 6754 800 12842 856
rect 13010 800 19098 856
rect 19266 800 21968 856
<< metal3 >>
rect 0 19048 800 19168
rect 21789 14696 22589 14816
rect 0 9800 800 9920
rect 21789 5448 22589 5568
<< obsm3 >>
rect 800 19248 21789 22337
rect 880 18968 21789 19248
rect 800 14896 21789 18968
rect 800 14616 21709 14896
rect 800 10000 21789 14616
rect 880 9720 21789 10000
rect 800 5648 21789 9720
rect 800 5368 21709 5648
rect 800 2143 21789 5368
<< metal4 >>
rect 4333 2128 4653 22352
rect 7721 2128 8041 22352
rect 11110 2128 11430 22352
rect 14499 2128 14819 22352
rect 17887 2128 18207 22352
<< obsm4 >>
rect 4733 2128 7641 22352
rect 8121 2128 11030 22352
rect 11510 2128 14419 22352
<< metal5 >>
rect 1104 18741 21436 19061
rect 1104 15387 21436 15707
rect 1104 12032 21436 12352
rect 1104 8677 21436 8997
rect 1104 5323 21436 5643
<< obsm5 >>
rect 1104 12672 21436 15067
rect 1104 9317 21436 11712
rect 1104 5963 21436 8357
<< labels >>
rlabel metal2 s 12898 0 12954 800 6 change[0]
port 1 nsew signal output
rlabel metal2 s 21914 23933 21970 24733 6 change[1]
port 2 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 choice[0]
port 3 nsew signal input
rlabel metal2 s 570 0 626 800 6 choice[1]
port 4 nsew signal input
rlabel metal3 s 21789 14696 22589 14816 6 choice[2]
port 5 nsew signal input
rlabel metal2 s 3330 23933 3386 24733 6 clk
port 6 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 coin[0]
port 7 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 coin[1]
port 8 nsew signal input
rlabel metal3 s 21789 5448 22589 5568 6 out[0]
port 9 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 out[1]
port 10 nsew signal output
rlabel metal2 s 15842 23933 15898 24733 6 out[2]
port 11 nsew signal output
rlabel metal2 s 9586 23933 9642 24733 6 reset
port 12 nsew signal input
rlabel metal4 s 17887 2128 18207 22352 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 11110 2128 11430 22352 6 VPWR
port 14 nsew power bidirectional
rlabel metal4 s 4333 2128 4653 22352 6 VPWR
port 15 nsew power bidirectional
rlabel metal5 s 1104 18741 21436 19061 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1104 12032 21436 12352 6 VPWR
port 17 nsew power bidirectional
rlabel metal5 s 1104 5323 21436 5643 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 14499 2128 14819 22352 6 VGND
port 19 nsew ground bidirectional
rlabel metal4 s 7721 2128 8041 22352 6 VGND
port 20 nsew ground bidirectional
rlabel metal5 s 1104 15387 21436 15707 6 VGND
port 21 nsew ground bidirectional
rlabel metal5 s 1104 8677 21436 8997 6 VGND
port 22 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22589 24733
string LEFview TRUE
<< end >>
