magic
tech sky130A
magscale 1 2
timestamp 1617727139
<< checkpaint >>
rect -3932 -3932 26521 28665
<< locali >>
rect 10057 9911 10091 10081
<< viali >>
rect 18337 22117 18371 22151
rect 18521 22049 18555 22083
rect 18613 21845 18647 21879
rect 18429 21641 18463 21675
rect 18318 21573 18352 21607
rect 18521 21505 18555 21539
rect 18613 21505 18647 21539
rect 9413 21437 9447 21471
rect 19717 21437 19751 21471
rect 19901 21437 19935 21471
rect 9229 21369 9263 21403
rect 9781 21369 9815 21403
rect 18153 21369 18187 21403
rect 19993 21301 20027 21335
rect 18981 21029 19015 21063
rect 19073 21029 19107 21063
rect 12449 20961 12483 20995
rect 12725 20961 12759 20995
rect 18889 20961 18923 20995
rect 12909 20893 12943 20927
rect 18705 20893 18739 20927
rect 19441 20893 19475 20927
rect 12541 20825 12575 20859
rect 13921 20349 13955 20383
rect 16865 20349 16899 20383
rect 20177 20349 20211 20383
rect 14013 20213 14047 20247
rect 16957 20213 16991 20247
rect 20269 20213 20303 20247
rect 2145 20009 2179 20043
rect 2513 19873 2547 19907
rect 2881 19873 2915 19907
rect 16405 19873 16439 19907
rect 16589 19873 16623 19907
rect 2605 19805 2639 19839
rect 2789 19805 2823 19839
rect 16681 19669 16715 19703
rect 1961 19261 1995 19295
rect 7481 19261 7515 19295
rect 7757 19261 7791 19295
rect 13369 19261 13403 19295
rect 13645 19261 13679 19295
rect 15025 19193 15059 19227
rect 2053 19125 2087 19159
rect 8861 19125 8895 19159
rect 17509 18853 17543 18887
rect 15853 18785 15887 18819
rect 16129 18717 16163 18751
rect 6837 18241 6871 18275
rect 7113 18173 7147 18207
rect 20085 18173 20119 18207
rect 7021 18105 7055 18139
rect 7573 18105 7607 18139
rect 20269 18037 20303 18071
rect 1409 17697 1443 17731
rect 1655 17697 1689 17731
rect 15945 17697 15979 17731
rect 16313 17697 16347 17731
rect 1869 17629 1903 17663
rect 15853 17629 15887 17663
rect 16405 17629 16439 17663
rect 1501 17561 1535 17595
rect 15393 17493 15427 17527
rect 4353 17085 4387 17119
rect 4721 17085 4755 17119
rect 4813 17085 4847 17119
rect 6837 17085 6871 17119
rect 3893 17017 3927 17051
rect 7021 16949 7055 16983
rect 16313 16677 16347 16711
rect 16865 16677 16899 16711
rect 13001 16609 13035 16643
rect 13093 16609 13127 16643
rect 16129 16609 16163 16643
rect 16405 16609 16439 16643
rect 2973 16201 3007 16235
rect 14289 16201 14323 16235
rect 7849 16065 7883 16099
rect 2881 15997 2915 16031
rect 7389 15997 7423 16031
rect 7665 15997 7699 16031
rect 14013 15997 14047 16031
rect 14105 15997 14139 16031
rect 6837 15929 6871 15963
rect 4813 15521 4847 15555
rect 15301 15521 15335 15555
rect 4905 15317 4939 15351
rect 15393 15317 15427 15351
rect 12725 14977 12759 15011
rect 13415 14977 13449 15011
rect 3525 14909 3559 14943
rect 3801 14909 3835 14943
rect 13277 14909 13311 14943
rect 13553 14909 13587 14943
rect 15301 14909 15335 14943
rect 15117 14841 15151 14875
rect 5089 14773 5123 14807
rect 15393 14773 15427 14807
rect 8493 14569 8527 14603
rect 4077 14433 4111 14467
rect 8677 14433 8711 14467
rect 9689 14433 9723 14467
rect 17969 14433 18003 14467
rect 18153 14433 18187 14467
rect 18337 14433 18371 14467
rect 4353 14365 4387 14399
rect 5733 14365 5767 14399
rect 17509 14365 17543 14399
rect 9873 14229 9907 14263
rect 17509 13481 17543 13515
rect 16865 13413 16899 13447
rect 17012 13277 17046 13311
rect 17233 13277 17267 13311
rect 17141 13209 17175 13243
rect 4813 12937 4847 12971
rect 14657 12937 14691 12971
rect 14197 12869 14231 12903
rect 3249 12801 3283 12835
rect 3525 12801 3559 12835
rect 14473 12733 14507 12767
rect 19625 12733 19659 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 14381 12665 14415 12699
rect 20085 12597 20119 12631
rect 10701 12257 10735 12291
rect 10977 12257 11011 12291
rect 12081 12053 12115 12087
rect 3525 11849 3559 11883
rect 16221 11849 16255 11883
rect 4261 11713 4295 11747
rect 3801 11645 3835 11679
rect 8677 11645 8711 11679
rect 12633 11645 12667 11679
rect 16129 11645 16163 11679
rect 3709 11577 3743 11611
rect 12449 11577 12483 11611
rect 12817 11577 12851 11611
rect 13185 11577 13219 11611
rect 15945 11577 15979 11611
rect 9965 11509 9999 11543
rect 12725 11509 12759 11543
rect 4997 11305 5031 11339
rect 6929 11305 6963 11339
rect 11069 11305 11103 11339
rect 4353 11237 4387 11271
rect 4583 11169 4617 11203
rect 6929 11169 6963 11203
rect 7573 11169 7607 11203
rect 7849 11169 7883 11203
rect 4721 11101 4755 11135
rect 9689 11101 9723 11135
rect 9965 11101 9999 11135
rect 4518 10965 4552 10999
rect 20085 10761 20119 10795
rect 9413 10625 9447 10659
rect 7113 10557 7147 10591
rect 7297 10557 7331 10591
rect 7665 10557 7699 10591
rect 8953 10557 8987 10591
rect 12909 10557 12943 10591
rect 13185 10557 13219 10591
rect 16313 10557 16347 10591
rect 19625 10557 19659 10591
rect 19809 10557 19843 10591
rect 19901 10557 19935 10591
rect 8677 10489 8711 10523
rect 8861 10489 8895 10523
rect 9045 10489 9079 10523
rect 16129 10489 16163 10523
rect 16681 10489 16715 10523
rect 14289 10421 14323 10455
rect 10149 10149 10183 10183
rect 16957 10149 16991 10183
rect 17325 10149 17359 10183
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 10057 10081 10091 10115
rect 10333 10081 10367 10115
rect 10701 10081 10735 10115
rect 16773 10081 16807 10115
rect 16865 10081 16899 10115
rect 18981 10081 19015 10115
rect 19349 10081 19383 10115
rect 2421 10013 2455 10047
rect 1777 9945 1811 9979
rect 16589 10013 16623 10047
rect 19625 10013 19659 10047
rect 18889 9945 18923 9979
rect 10057 9877 10091 9911
rect 9045 9469 9079 9503
rect 19993 9469 20027 9503
rect 8861 9333 8895 9367
rect 20177 9333 20211 9367
rect 3065 9061 3099 9095
rect 13829 9061 13863 9095
rect 13921 9061 13955 9095
rect 14381 9061 14415 9095
rect 1409 8993 1443 9027
rect 9781 8993 9815 9027
rect 9873 8993 9907 9027
rect 11161 8993 11195 9027
rect 13997 8993 14031 9027
rect 1685 8925 1719 8959
rect 11253 8925 11287 8959
rect 13645 8925 13679 8959
rect 10057 8789 10091 8823
rect 3617 8585 3651 8619
rect 8401 8517 8435 8551
rect 15945 8449 15979 8483
rect 3525 8381 3559 8415
rect 7021 8381 7055 8415
rect 7297 8381 7331 8415
rect 15209 8381 15243 8415
rect 15393 8381 15427 8415
rect 15485 8381 15519 8415
rect 15577 8313 15611 8347
rect 17325 8041 17359 8075
rect 4629 7973 4663 8007
rect 2421 7905 2455 7939
rect 4077 7905 4111 7939
rect 4169 7905 4203 7939
rect 16865 7905 16899 7939
rect 17141 7905 17175 7939
rect 2513 7769 2547 7803
rect 16957 7769 16991 7803
rect 15485 7497 15519 7531
rect 4629 7361 4663 7395
rect 10149 7361 10183 7395
rect 1409 7293 1443 7327
rect 3157 7293 3191 7327
rect 3341 7293 3375 7327
rect 3525 7293 3559 7327
rect 3801 7293 3835 7327
rect 4054 7293 4088 7327
rect 9781 7293 9815 7327
rect 15393 7293 15427 7327
rect 9597 7225 9631 7259
rect 15209 7225 15243 7259
rect 1593 7157 1627 7191
rect 2789 6885 2823 6919
rect 2053 6817 2087 6851
rect 2329 6817 2363 6851
rect 10241 6817 10275 6851
rect 10333 6817 10367 6851
rect 15301 6817 15335 6851
rect 15448 6817 15482 6851
rect 19441 6817 19475 6851
rect 19625 6817 19659 6851
rect 2145 6749 2179 6783
rect 7021 6749 7055 6783
rect 7297 6749 7331 6783
rect 15669 6749 15703 6783
rect 15577 6681 15611 6715
rect 8401 6613 8435 6647
rect 15761 6613 15795 6647
rect 19717 6613 19751 6647
rect 2605 6341 2639 6375
rect 2789 6205 2823 6239
rect 2973 6205 3007 6239
rect 3157 6205 3191 6239
rect 11529 5865 11563 5899
rect 2605 5797 2639 5831
rect 10885 5797 10919 5831
rect 2717 5729 2751 5763
rect 3157 5729 3191 5763
rect 11032 5729 11066 5763
rect 11253 5661 11287 5695
rect 2421 5593 2455 5627
rect 11161 5593 11195 5627
rect 1501 4777 1535 4811
rect 6377 4777 6411 4811
rect 17325 4777 17359 4811
rect 1401 4641 1435 4675
rect 6469 4641 6503 4675
rect 6837 4641 6871 4675
rect 7113 4641 7147 4675
rect 16221 4641 16255 4675
rect 15945 4573 15979 4607
rect 7757 4233 7791 4267
rect 3157 4097 3191 4131
rect 3893 4097 3927 4131
rect 8493 4097 8527 4131
rect 3801 4029 3835 4063
rect 4169 4029 4203 4063
rect 4353 4029 4387 4063
rect 7941 4029 7975 4063
rect 8033 4029 8067 4063
rect 12541 4029 12575 4063
rect 12725 4029 12759 4063
rect 12817 4029 12851 4063
rect 13277 3961 13311 3995
rect 10793 3689 10827 3723
rect 10701 3553 10735 3587
rect 4445 3009 4479 3043
rect 5181 3009 5215 3043
rect 4721 2941 4755 2975
rect 20085 2941 20119 2975
rect 4813 2873 4847 2907
rect 4629 2805 4663 2839
rect 20269 2805 20303 2839
rect 10517 2533 10551 2567
rect 6929 2465 6963 2499
rect 7021 2465 7055 2499
rect 11069 2465 11103 2499
rect 11345 2465 11379 2499
rect 11529 2465 11563 2499
rect 7481 2397 7515 2431
<< metal1 >>
rect 1104 22330 21436 22352
rect 1104 22278 7759 22330
rect 7811 22278 7823 22330
rect 7875 22278 7887 22330
rect 7939 22278 7951 22330
rect 8003 22278 14536 22330
rect 14588 22278 14600 22330
rect 14652 22278 14664 22330
rect 14716 22278 14728 22330
rect 14780 22278 21436 22330
rect 1104 22256 21436 22278
rect 8570 22108 8576 22160
rect 8628 22148 8634 22160
rect 18325 22151 18383 22157
rect 18325 22148 18337 22151
rect 8628 22120 18337 22148
rect 8628 22108 8634 22120
rect 18325 22117 18337 22120
rect 18371 22117 18383 22151
rect 18325 22111 18383 22117
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 18509 22083 18567 22089
rect 18509 22080 18521 22083
rect 15344 22052 18521 22080
rect 15344 22040 15350 22052
rect 18509 22049 18521 22052
rect 18555 22049 18567 22083
rect 18509 22043 18567 22049
rect 7374 21904 7380 21956
rect 7432 21944 7438 21956
rect 19702 21944 19708 21956
rect 7432 21916 19708 21944
rect 7432 21904 7438 21916
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 13504 21848 18613 21876
rect 13504 21836 13510 21848
rect 18601 21845 18613 21848
rect 18647 21845 18659 21879
rect 18601 21839 18659 21845
rect 1104 21786 21436 21808
rect 1104 21734 4370 21786
rect 4422 21734 4434 21786
rect 4486 21734 4498 21786
rect 4550 21734 4562 21786
rect 4614 21734 11148 21786
rect 11200 21734 11212 21786
rect 11264 21734 11276 21786
rect 11328 21734 11340 21786
rect 11392 21734 17925 21786
rect 17977 21734 17989 21786
rect 18041 21734 18053 21786
rect 18105 21734 18117 21786
rect 18169 21734 21436 21786
rect 1104 21712 21436 21734
rect 18417 21675 18475 21681
rect 18417 21672 18429 21675
rect 14016 21644 18429 21672
rect 12066 21564 12072 21616
rect 12124 21604 12130 21616
rect 14016 21604 14044 21644
rect 18417 21641 18429 21644
rect 18463 21641 18475 21675
rect 18417 21635 18475 21641
rect 12124 21576 14044 21604
rect 18306 21607 18364 21613
rect 12124 21564 12130 21576
rect 18306 21573 18318 21607
rect 18352 21604 18364 21607
rect 18966 21604 18972 21616
rect 18352 21576 18972 21604
rect 18352 21573 18364 21576
rect 18306 21567 18364 21573
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 18509 21539 18567 21545
rect 18509 21536 18521 21539
rect 12032 21508 18521 21536
rect 12032 21496 12038 21508
rect 18509 21505 18521 21508
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 18601 21539 18659 21545
rect 18601 21505 18613 21539
rect 18647 21505 18659 21539
rect 18601 21499 18659 21505
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 13170 21468 13176 21480
rect 9447 21440 13176 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 18616 21468 18644 21499
rect 19702 21468 19708 21480
rect 17000 21440 18644 21468
rect 19663 21440 19708 21468
rect 17000 21428 17006 21440
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 19886 21468 19892 21480
rect 19847 21440 19892 21468
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 9214 21400 9220 21412
rect 9175 21372 9220 21400
rect 9214 21360 9220 21372
rect 9272 21360 9278 21412
rect 9769 21403 9827 21409
rect 9769 21369 9781 21403
rect 9815 21400 9827 21403
rect 16298 21400 16304 21412
rect 9815 21372 16304 21400
rect 9815 21369 9827 21372
rect 9769 21363 9827 21369
rect 16298 21360 16304 21372
rect 16356 21400 16362 21412
rect 18141 21403 18199 21409
rect 18141 21400 18153 21403
rect 16356 21372 18153 21400
rect 16356 21360 16362 21372
rect 18141 21369 18153 21372
rect 18187 21369 18199 21403
rect 18141 21363 18199 21369
rect 18248 21372 20024 21400
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 18248 21332 18276 21372
rect 19996 21341 20024 21372
rect 16632 21304 18276 21332
rect 19981 21335 20039 21341
rect 16632 21292 16638 21304
rect 19981 21301 19993 21335
rect 20027 21301 20039 21335
rect 19981 21295 20039 21301
rect 1104 21242 21436 21264
rect 1104 21190 7759 21242
rect 7811 21190 7823 21242
rect 7875 21190 7887 21242
rect 7939 21190 7951 21242
rect 8003 21190 14536 21242
rect 14588 21190 14600 21242
rect 14652 21190 14664 21242
rect 14716 21190 14728 21242
rect 14780 21190 21436 21242
rect 1104 21168 21436 21190
rect 17586 21088 17592 21140
rect 17644 21128 17650 21140
rect 19886 21128 19892 21140
rect 17644 21100 19892 21128
rect 17644 21088 17650 21100
rect 19886 21088 19892 21100
rect 19944 21088 19950 21140
rect 16758 21020 16764 21072
rect 16816 21060 16822 21072
rect 18969 21063 19027 21069
rect 18969 21060 18981 21063
rect 16816 21032 18981 21060
rect 16816 21020 16822 21032
rect 18969 21029 18981 21032
rect 19015 21029 19027 21063
rect 18969 21023 19027 21029
rect 19061 21063 19119 21069
rect 19061 21029 19073 21063
rect 19107 21060 19119 21063
rect 20254 21060 20260 21072
rect 19107 21032 20260 21060
rect 19107 21029 19119 21032
rect 19061 21023 19119 21029
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 12437 20995 12495 21001
rect 12437 20992 12449 20995
rect 6420 20964 12449 20992
rect 6420 20952 6426 20964
rect 12437 20961 12449 20964
rect 12483 20961 12495 20995
rect 12710 20992 12716 21004
rect 12671 20964 12716 20992
rect 12437 20955 12495 20961
rect 12710 20952 12716 20964
rect 12768 20952 12774 21004
rect 16390 20952 16396 21004
rect 16448 20992 16454 21004
rect 18877 20995 18935 21001
rect 18877 20992 18889 20995
rect 16448 20964 18889 20992
rect 16448 20952 16454 20964
rect 18877 20961 18889 20964
rect 18923 20961 18935 20995
rect 18877 20955 18935 20961
rect 10686 20884 10692 20936
rect 10744 20924 10750 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 10744 20896 12909 20924
rect 10744 20884 10750 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 16666 20884 16672 20936
rect 16724 20924 16730 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 16724 20896 18705 20924
rect 16724 20884 16730 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 8294 20816 8300 20868
rect 8352 20856 8358 20868
rect 12529 20859 12587 20865
rect 12529 20856 12541 20859
rect 8352 20828 12541 20856
rect 8352 20816 8358 20828
rect 12529 20825 12541 20828
rect 12575 20825 12587 20859
rect 12529 20819 12587 20825
rect 17402 20816 17408 20868
rect 17460 20856 17466 20868
rect 19444 20856 19472 20887
rect 17460 20828 19472 20856
rect 17460 20816 17466 20828
rect 1104 20698 21436 20720
rect 1104 20646 4370 20698
rect 4422 20646 4434 20698
rect 4486 20646 4498 20698
rect 4550 20646 4562 20698
rect 4614 20646 11148 20698
rect 11200 20646 11212 20698
rect 11264 20646 11276 20698
rect 11328 20646 11340 20698
rect 11392 20646 17925 20698
rect 17977 20646 17989 20698
rect 18041 20646 18053 20698
rect 18105 20646 18117 20698
rect 18169 20646 21436 20698
rect 1104 20624 21436 20646
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 12158 20584 12164 20596
rect 9640 20556 12164 20584
rect 9640 20544 9646 20556
rect 12158 20544 12164 20556
rect 12216 20584 12222 20596
rect 12710 20584 12716 20596
rect 12216 20556 12716 20584
rect 12216 20544 12222 20556
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12768 20420 20208 20448
rect 12768 20408 12774 20420
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20380 13967 20383
rect 14826 20380 14832 20392
rect 13955 20352 14832 20380
rect 13955 20349 13967 20352
rect 13909 20343 13967 20349
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 16853 20383 16911 20389
rect 16853 20349 16865 20383
rect 16899 20380 16911 20383
rect 17494 20380 17500 20392
rect 16899 20352 17500 20380
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 20180 20389 20208 20420
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 8386 20272 8392 20324
rect 8444 20312 8450 20324
rect 15838 20312 15844 20324
rect 8444 20284 15844 20312
rect 8444 20272 8450 20284
rect 15838 20272 15844 20284
rect 15896 20272 15902 20324
rect 14001 20247 14059 20253
rect 14001 20213 14013 20247
rect 14047 20244 14059 20247
rect 15102 20244 15108 20256
rect 14047 20216 15108 20244
rect 14047 20213 14059 20216
rect 14001 20207 14059 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 16945 20247 17003 20253
rect 16945 20213 16957 20247
rect 16991 20244 17003 20247
rect 17034 20244 17040 20256
rect 16991 20216 17040 20244
rect 16991 20213 17003 20216
rect 16945 20207 17003 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 20257 20247 20315 20253
rect 20257 20244 20269 20247
rect 19392 20216 20269 20244
rect 19392 20204 19398 20216
rect 20257 20213 20269 20216
rect 20303 20213 20315 20247
rect 20257 20207 20315 20213
rect 1104 20154 21436 20176
rect 1104 20102 7759 20154
rect 7811 20102 7823 20154
rect 7875 20102 7887 20154
rect 7939 20102 7951 20154
rect 8003 20102 14536 20154
rect 14588 20102 14600 20154
rect 14652 20102 14664 20154
rect 14716 20102 14728 20154
rect 14780 20102 21436 20154
rect 1104 20080 21436 20102
rect 2133 20043 2191 20049
rect 2133 20009 2145 20043
rect 2179 20040 2191 20043
rect 10134 20040 10140 20052
rect 2179 20012 10140 20040
rect 2179 20009 2191 20012
rect 2133 20003 2191 20009
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 2958 19972 2964 19984
rect 2516 19944 2964 19972
rect 2516 19913 2544 19944
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 21910 19972 21916 19984
rect 8904 19944 21916 19972
rect 8904 19932 8910 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 11514 19904 11520 19916
rect 2915 19876 11520 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 16390 19904 16396 19916
rect 16351 19876 16396 19904
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 16577 19907 16635 19913
rect 16577 19873 16589 19907
rect 16623 19904 16635 19907
rect 16666 19904 16672 19916
rect 16623 19876 16672 19904
rect 16623 19873 16635 19876
rect 16577 19867 16635 19873
rect 16666 19864 16672 19876
rect 16724 19864 16730 19916
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19805 2651 19839
rect 2593 19799 2651 19805
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 11790 19836 11796 19848
rect 2823 19808 11796 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 2608 19768 2636 19799
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 17586 19836 17592 19848
rect 11992 19808 17592 19836
rect 11992 19768 12020 19808
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 2608 19740 12020 19768
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 16669 19703 16727 19709
rect 16669 19700 16681 19703
rect 15068 19672 16681 19700
rect 15068 19660 15074 19672
rect 16669 19669 16681 19672
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 1104 19610 21436 19632
rect 1104 19558 4370 19610
rect 4422 19558 4434 19610
rect 4486 19558 4498 19610
rect 4550 19558 4562 19610
rect 4614 19558 11148 19610
rect 11200 19558 11212 19610
rect 11264 19558 11276 19610
rect 11328 19558 11340 19610
rect 11392 19558 17925 19610
rect 17977 19558 17989 19610
rect 18041 19558 18053 19610
rect 18105 19558 18117 19610
rect 18169 19558 21436 19610
rect 1104 19536 21436 19558
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 8662 19360 8668 19372
rect 3384 19332 8668 19360
rect 3384 19320 3390 19332
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19292 7803 19295
rect 8110 19292 8116 19304
rect 7791 19264 8116 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 7374 19156 7380 19168
rect 2087 19128 7380 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 7484 19156 7512 19255
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 13354 19292 13360 19304
rect 8404 19264 13360 19292
rect 8404 19156 8432 19264
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13630 19292 13636 19304
rect 13591 19264 13636 19292
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 15013 19227 15071 19233
rect 15013 19193 15025 19227
rect 15059 19224 15071 19227
rect 16482 19224 16488 19236
rect 15059 19196 16488 19224
rect 15059 19193 15071 19196
rect 15013 19187 15071 19193
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 8478 19156 8484 19168
rect 7484 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 1104 19066 21436 19088
rect 1104 19014 7759 19066
rect 7811 19014 7823 19066
rect 7875 19014 7887 19066
rect 7939 19014 7951 19066
rect 8003 19014 14536 19066
rect 14588 19014 14600 19066
rect 14652 19014 14664 19066
rect 14716 19014 14728 19066
rect 14780 19014 21436 19066
rect 1104 18992 21436 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 17310 18952 17316 18964
rect 2004 18924 17316 18952
rect 2004 18912 2010 18924
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 17218 18844 17224 18896
rect 17276 18884 17282 18896
rect 17497 18887 17555 18893
rect 17497 18884 17509 18887
rect 17276 18856 17509 18884
rect 17276 18844 17282 18856
rect 17497 18853 17509 18856
rect 17543 18884 17555 18887
rect 17586 18884 17592 18896
rect 17543 18856 17592 18884
rect 17543 18853 17555 18856
rect 17497 18847 17555 18853
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 13412 18788 15853 18816
rect 13412 18776 13418 18788
rect 15841 18785 15853 18788
rect 15887 18785 15899 18819
rect 15841 18779 15899 18785
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16850 18748 16856 18760
rect 16163 18720 16856 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 1104 18522 21436 18544
rect 1104 18470 4370 18522
rect 4422 18470 4434 18522
rect 4486 18470 4498 18522
rect 4550 18470 4562 18522
rect 4614 18470 11148 18522
rect 11200 18470 11212 18522
rect 11264 18470 11276 18522
rect 11328 18470 11340 18522
rect 11392 18470 17925 18522
rect 17977 18470 17989 18522
rect 18041 18470 18053 18522
rect 18105 18470 18117 18522
rect 18169 18470 21436 18522
rect 1104 18448 21436 18470
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 11698 18272 11704 18284
rect 6871 18244 11704 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 7101 18207 7159 18213
rect 7101 18204 7113 18207
rect 6932 18176 7113 18204
rect 3602 18096 3608 18148
rect 3660 18136 3666 18148
rect 6932 18136 6960 18176
rect 7101 18173 7113 18176
rect 7147 18173 7159 18207
rect 7101 18167 7159 18173
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 18966 18204 18972 18216
rect 13320 18176 18972 18204
rect 13320 18164 13326 18176
rect 18966 18164 18972 18176
rect 19024 18204 19030 18216
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19024 18176 20085 18204
rect 19024 18164 19030 18176
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 20073 18167 20131 18173
rect 3660 18108 6960 18136
rect 7009 18139 7067 18145
rect 3660 18096 3666 18108
rect 7009 18105 7021 18139
rect 7055 18105 7067 18139
rect 7558 18136 7564 18148
rect 7519 18108 7564 18136
rect 7009 18099 7067 18105
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 7024 18068 7052 18099
rect 7558 18096 7564 18108
rect 7616 18096 7622 18148
rect 20254 18068 20260 18080
rect 6972 18040 7052 18068
rect 20215 18040 20260 18068
rect 6972 18028 6978 18040
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 1104 17978 21436 18000
rect 1104 17926 7759 17978
rect 7811 17926 7823 17978
rect 7875 17926 7887 17978
rect 7939 17926 7951 17978
rect 8003 17926 14536 17978
rect 14588 17926 14600 17978
rect 14652 17926 14664 17978
rect 14716 17926 14728 17978
rect 14780 17926 21436 17978
rect 1104 17904 21436 17926
rect 12158 17796 12164 17808
rect 1688 17768 12164 17796
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1688 17737 1716 17768
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 14366 17756 14372 17808
rect 14424 17796 14430 17808
rect 14424 17768 16344 17796
rect 14424 17756 14430 17768
rect 1643 17731 1716 17737
rect 1643 17697 1655 17731
rect 1689 17700 1716 17731
rect 1689 17697 1701 17700
rect 1643 17691 1701 17697
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 16316 17737 16344 17768
rect 15933 17731 15991 17737
rect 15933 17728 15945 17731
rect 10468 17700 15945 17728
rect 10468 17688 10474 17700
rect 15933 17697 15945 17700
rect 15979 17697 15991 17731
rect 15933 17691 15991 17697
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 1854 17660 1860 17672
rect 1815 17632 1860 17660
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 11664 17632 15853 17660
rect 11664 17620 11670 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 1489 17595 1547 17601
rect 1489 17561 1501 17595
rect 1535 17592 1547 17595
rect 2682 17592 2688 17604
rect 1535 17564 2688 17592
rect 1535 17561 1547 17564
rect 1489 17555 1547 17561
rect 2682 17552 2688 17564
rect 2740 17552 2746 17604
rect 15654 17552 15660 17604
rect 15712 17592 15718 17604
rect 16408 17592 16436 17623
rect 15712 17564 16436 17592
rect 15712 17552 15718 17564
rect 15378 17524 15384 17536
rect 15339 17496 15384 17524
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 1104 17434 21436 17456
rect 1104 17382 4370 17434
rect 4422 17382 4434 17434
rect 4486 17382 4498 17434
rect 4550 17382 4562 17434
rect 4614 17382 11148 17434
rect 11200 17382 11212 17434
rect 11264 17382 11276 17434
rect 11328 17382 11340 17434
rect 11392 17382 17925 17434
rect 17977 17382 17989 17434
rect 18041 17382 18053 17434
rect 18105 17382 18117 17434
rect 18169 17382 21436 17434
rect 1104 17360 21436 17382
rect 17034 17320 17040 17332
rect 4356 17292 17040 17320
rect 4356 17125 4384 17292
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 5350 17184 5356 17196
rect 4724 17156 5356 17184
rect 4724 17125 4752 17156
rect 5350 17144 5356 17156
rect 5408 17184 5414 17196
rect 13078 17184 13084 17196
rect 5408 17156 13084 17184
rect 5408 17144 5414 17156
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 5258 17116 5264 17128
rect 4847 17088 5264 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6788 17088 6837 17116
rect 6788 17076 6794 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 3786 17008 3792 17060
rect 3844 17048 3850 17060
rect 3881 17051 3939 17057
rect 3881 17048 3893 17051
rect 3844 17020 3893 17048
rect 3844 17008 3850 17020
rect 3881 17017 3893 17020
rect 3927 17048 3939 17051
rect 15286 17048 15292 17060
rect 3927 17020 15292 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 7009 16983 7067 16989
rect 7009 16949 7021 16983
rect 7055 16980 7067 16983
rect 9490 16980 9496 16992
rect 7055 16952 9496 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 9490 16940 9496 16952
rect 9548 16980 9554 16992
rect 16390 16980 16396 16992
rect 9548 16952 16396 16980
rect 9548 16940 9554 16952
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 1104 16890 21436 16912
rect 1104 16838 7759 16890
rect 7811 16838 7823 16890
rect 7875 16838 7887 16890
rect 7939 16838 7951 16890
rect 8003 16838 14536 16890
rect 14588 16838 14600 16890
rect 14652 16838 14664 16890
rect 14716 16838 14728 16890
rect 14780 16838 21436 16890
rect 1104 16816 21436 16838
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14056 16748 16252 16776
rect 14056 16736 14062 16748
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 11756 16680 16160 16708
rect 11756 16668 11762 16680
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 12986 16640 12992 16652
rect 3016 16612 12992 16640
rect 3016 16600 3022 16612
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 16132 16649 16160 16680
rect 16117 16643 16175 16649
rect 13136 16612 13181 16640
rect 13136 16600 13142 16612
rect 16117 16609 16129 16643
rect 16163 16609 16175 16643
rect 16224 16640 16252 16748
rect 16301 16711 16359 16717
rect 16301 16677 16313 16711
rect 16347 16708 16359 16711
rect 16574 16708 16580 16720
rect 16347 16680 16580 16708
rect 16347 16677 16359 16680
rect 16301 16671 16359 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 16850 16708 16856 16720
rect 16811 16680 16856 16708
rect 16850 16668 16856 16680
rect 16908 16668 16914 16720
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 16224 16612 16405 16640
rect 16117 16603 16175 16609
rect 16393 16609 16405 16612
rect 16439 16609 16451 16643
rect 16393 16603 16451 16609
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 16758 16572 16764 16584
rect 16632 16544 16764 16572
rect 16632 16532 16638 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 1104 16346 21436 16368
rect 1104 16294 4370 16346
rect 4422 16294 4434 16346
rect 4486 16294 4498 16346
rect 4550 16294 4562 16346
rect 4614 16294 11148 16346
rect 11200 16294 11212 16346
rect 11264 16294 11276 16346
rect 11328 16294 11340 16346
rect 11392 16294 17925 16346
rect 17977 16294 17989 16346
rect 18041 16294 18053 16346
rect 18105 16294 18117 16346
rect 18169 16294 21436 16346
rect 1104 16272 21436 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 6730 16232 6736 16244
rect 3007 16204 6736 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 14274 16232 14280 16244
rect 14235 16204 14280 16232
rect 14274 16192 14280 16204
rect 14332 16192 14338 16244
rect 7837 16099 7895 16105
rect 7837 16096 7849 16099
rect 5276 16068 7849 16096
rect 2866 16028 2872 16040
rect 2827 16000 2872 16028
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 2406 15920 2412 15972
rect 2464 15960 2470 15972
rect 2682 15960 2688 15972
rect 2464 15932 2688 15960
rect 2464 15920 2470 15932
rect 2682 15920 2688 15932
rect 2740 15960 2746 15972
rect 5276 15960 5304 16068
rect 7837 16065 7849 16068
rect 7883 16065 7895 16099
rect 7837 16059 7895 16065
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7374 16028 7380 16040
rect 7156 16000 7380 16028
rect 7156 15988 7162 16000
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 7650 16028 7656 16040
rect 7611 16000 7656 16028
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14182 16028 14188 16040
rect 14139 16000 14188 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 2740 15932 5304 15960
rect 6825 15963 6883 15969
rect 2740 15920 2746 15932
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 8294 15960 8300 15972
rect 6871 15932 8300 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 6730 15852 6736 15904
rect 6788 15892 6794 15904
rect 9950 15892 9956 15904
rect 6788 15864 9956 15892
rect 6788 15852 6794 15864
rect 9950 15852 9956 15864
rect 10008 15892 10014 15904
rect 14016 15892 14044 15991
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 10008 15864 14044 15892
rect 10008 15852 10014 15864
rect 1104 15802 21436 15824
rect 1104 15750 7759 15802
rect 7811 15750 7823 15802
rect 7875 15750 7887 15802
rect 7939 15750 7951 15802
rect 8003 15750 14536 15802
rect 14588 15750 14600 15802
rect 14652 15750 14664 15802
rect 14716 15750 14728 15802
rect 14780 15750 21436 15802
rect 1104 15728 21436 15750
rect 2866 15580 2872 15632
rect 2924 15620 2930 15632
rect 13722 15620 13728 15632
rect 2924 15592 13728 15620
rect 2924 15580 2930 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5074 15552 5080 15564
rect 4847 15524 5080 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 4890 15348 4896 15360
rect 4851 15320 4896 15348
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15381 15351 15439 15357
rect 15381 15348 15393 15351
rect 15252 15320 15393 15348
rect 15252 15308 15258 15320
rect 15381 15317 15393 15320
rect 15427 15317 15439 15351
rect 15381 15311 15439 15317
rect 1104 15258 21436 15280
rect 1104 15206 4370 15258
rect 4422 15206 4434 15258
rect 4486 15206 4498 15258
rect 4550 15206 4562 15258
rect 4614 15206 11148 15258
rect 11200 15206 11212 15258
rect 11264 15206 11276 15258
rect 11328 15206 11340 15258
rect 11392 15206 17925 15258
rect 17977 15206 17989 15258
rect 18041 15206 18053 15258
rect 18105 15206 18117 15258
rect 18169 15206 21436 15258
rect 1104 15184 21436 15206
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 12713 15011 12771 15017
rect 12713 15008 12725 15011
rect 11572 14980 12725 15008
rect 11572 14968 11578 14980
rect 12713 14977 12725 14980
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 13170 14968 13176 15020
rect 13228 15008 13234 15020
rect 13403 15011 13461 15017
rect 13403 15008 13415 15011
rect 13228 14980 13415 15008
rect 13228 14968 13234 14980
rect 13403 14977 13415 14980
rect 13449 14977 13461 15011
rect 14274 15008 14280 15020
rect 13403 14971 13461 14977
rect 13556 14980 14280 15008
rect 3510 14940 3516 14952
rect 3471 14912 3516 14940
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4246 14940 4252 14952
rect 3835 14912 4252 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 13556 14949 13584 14980
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13280 14872 13308 14903
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 13964 14912 15301 14940
rect 13964 14900 13970 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 14090 14872 14096 14884
rect 13280 14844 14096 14872
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 15838 14872 15844 14884
rect 15151 14844 15844 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 12434 14804 12440 14816
rect 5123 14776 12440 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 15381 14807 15439 14813
rect 15381 14804 15393 14807
rect 13872 14776 15393 14804
rect 13872 14764 13878 14776
rect 15381 14773 15393 14776
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 1104 14714 21436 14736
rect 1104 14662 7759 14714
rect 7811 14662 7823 14714
rect 7875 14662 7887 14714
rect 7939 14662 7951 14714
rect 8003 14662 14536 14714
rect 14588 14662 14600 14714
rect 14652 14662 14664 14714
rect 14716 14662 14728 14714
rect 14780 14662 21436 14714
rect 1104 14640 21436 14662
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3510 14600 3516 14612
rect 3292 14572 3516 14600
rect 3292 14560 3298 14572
rect 3510 14560 3516 14572
rect 3568 14600 3574 14612
rect 8478 14600 8484 14612
rect 3568 14572 8484 14600
rect 3568 14560 3574 14572
rect 4080 14473 4108 14572
rect 8478 14560 8484 14572
rect 8536 14600 8542 14612
rect 9030 14600 9036 14612
rect 8536 14572 9036 14600
rect 8536 14560 8542 14572
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 10042 14600 10048 14612
rect 9692 14572 10048 14600
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 9582 14464 9588 14476
rect 8711 14436 9588 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 9692 14473 9720 14572
rect 10042 14560 10048 14572
rect 10100 14600 10106 14612
rect 19334 14600 19340 14612
rect 10100 14572 19340 14600
rect 10100 14560 10106 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 13136 14504 18184 14532
rect 13136 14492 13142 14504
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 18156 14473 18184 14504
rect 17957 14467 18015 14473
rect 17957 14464 17969 14467
rect 17092 14436 17969 14464
rect 17092 14424 17098 14436
rect 17957 14433 17969 14436
rect 18003 14433 18015 14467
rect 17957 14427 18015 14433
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14433 18199 14467
rect 18141 14427 18199 14433
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18288 14436 18337 14464
rect 18288 14424 18294 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 5166 14396 5172 14408
rect 4387 14368 5172 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14396 5779 14399
rect 13262 14396 13268 14408
rect 5767 14368 13268 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 5736 14260 5764 14359
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17368 14368 17509 14396
rect 17368 14356 17374 14368
rect 17497 14365 17509 14368
rect 17543 14396 17555 14399
rect 17770 14396 17776 14408
rect 17543 14368 17776 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 4120 14232 5764 14260
rect 4120 14220 4126 14232
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9732 14232 9873 14260
rect 9732 14220 9738 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 9861 14223 9919 14229
rect 1104 14170 21436 14192
rect 1104 14118 4370 14170
rect 4422 14118 4434 14170
rect 4486 14118 4498 14170
rect 4550 14118 4562 14170
rect 4614 14118 11148 14170
rect 11200 14118 11212 14170
rect 11264 14118 11276 14170
rect 11328 14118 11340 14170
rect 11392 14118 17925 14170
rect 17977 14118 17989 14170
rect 18041 14118 18053 14170
rect 18105 14118 18117 14170
rect 18169 14118 21436 14170
rect 1104 14096 21436 14118
rect 1104 13626 21436 13648
rect 1104 13574 7759 13626
rect 7811 13574 7823 13626
rect 7875 13574 7887 13626
rect 7939 13574 7951 13626
rect 8003 13574 14536 13626
rect 14588 13574 14600 13626
rect 14652 13574 14664 13626
rect 14716 13574 14728 13626
rect 14780 13574 21436 13626
rect 1104 13552 21436 13574
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17494 13512 17500 13524
rect 17368 13484 17500 13512
rect 17368 13472 17374 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 16853 13447 16911 13453
rect 16853 13444 16865 13447
rect 16816 13416 16865 13444
rect 16816 13404 16822 13416
rect 16853 13413 16865 13416
rect 16899 13444 16911 13447
rect 16942 13444 16948 13456
rect 16899 13416 16948 13444
rect 16899 13413 16911 13416
rect 16853 13407 16911 13413
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 6972 13348 14688 13376
rect 6972 13336 6978 13348
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 13630 13308 13636 13320
rect 3936 13280 13636 13308
rect 3936 13268 3942 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14660 13308 14688 13348
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 17126 13376 17132 13388
rect 16540 13348 17132 13376
rect 16540 13336 16546 13348
rect 17126 13336 17132 13348
rect 17184 13376 17190 13388
rect 17184 13348 17264 13376
rect 17184 13336 17190 13348
rect 17236 13317 17264 13348
rect 17000 13311 17058 13317
rect 17000 13308 17012 13311
rect 14660 13280 17012 13308
rect 17000 13277 17012 13280
rect 17046 13277 17058 13311
rect 17000 13271 17058 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 3050 13200 3056 13252
rect 3108 13240 3114 13252
rect 17129 13243 17187 13249
rect 17129 13240 17141 13243
rect 3108 13212 17141 13240
rect 3108 13200 3114 13212
rect 17129 13209 17141 13212
rect 17175 13209 17187 13243
rect 17129 13203 17187 13209
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 15378 13172 15384 13184
rect 13504 13144 15384 13172
rect 13504 13132 13510 13144
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 1104 13082 21436 13104
rect 1104 13030 4370 13082
rect 4422 13030 4434 13082
rect 4486 13030 4498 13082
rect 4550 13030 4562 13082
rect 4614 13030 11148 13082
rect 11200 13030 11212 13082
rect 11264 13030 11276 13082
rect 11328 13030 11340 13082
rect 11392 13030 17925 13082
rect 17977 13030 17989 13082
rect 18041 13030 18053 13082
rect 18105 13030 18117 13082
rect 18169 13030 21436 13082
rect 1104 13008 21436 13030
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 3476 12940 4813 12968
rect 3476 12928 3482 12940
rect 4801 12937 4813 12940
rect 4847 12968 4859 12971
rect 6914 12968 6920 12980
rect 4847 12940 6920 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 13688 12940 14657 12968
rect 13688 12928 13694 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 14645 12931 14703 12937
rect 13446 12900 13452 12912
rect 10336 12872 13452 12900
rect 3234 12832 3240 12844
rect 3195 12804 3240 12832
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 10336 12832 10364 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 14185 12903 14243 12909
rect 14185 12900 14197 12903
rect 14148 12872 14197 12900
rect 14148 12860 14154 12872
rect 14185 12869 14197 12872
rect 14231 12900 14243 12903
rect 14918 12900 14924 12912
rect 14231 12872 14924 12900
rect 14231 12869 14243 12872
rect 14185 12863 14243 12869
rect 14918 12860 14924 12872
rect 14976 12860 14982 12912
rect 3559 12804 10364 12832
rect 13464 12804 14412 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 13464 12764 13492 12804
rect 14274 12764 14280 12776
rect 11848 12736 13492 12764
rect 14016 12736 14280 12764
rect 11848 12724 11854 12736
rect 14016 12640 14044 12736
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14384 12764 14412 12804
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 19300 12804 19932 12832
rect 19300 12792 19306 12804
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 14384 12736 14473 12764
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 19904 12773 19932 12804
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 15160 12736 19625 12764
rect 15160 12724 15166 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 14366 12696 14372 12708
rect 14279 12668 14372 12696
rect 14366 12656 14372 12668
rect 14424 12696 14430 12708
rect 15010 12696 15016 12708
rect 14424 12668 15016 12696
rect 14424 12656 14430 12668
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 11698 12628 11704 12640
rect 9180 12600 11704 12628
rect 9180 12588 9186 12600
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 13998 12588 14004 12640
rect 14056 12588 14062 12640
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 19720 12628 19748 12727
rect 20070 12628 20076 12640
rect 14332 12600 19748 12628
rect 20031 12600 20076 12628
rect 14332 12588 14338 12600
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 1104 12538 21436 12560
rect 1104 12486 7759 12538
rect 7811 12486 7823 12538
rect 7875 12486 7887 12538
rect 7939 12486 7951 12538
rect 8003 12486 14536 12538
rect 14588 12486 14600 12538
rect 14652 12486 14664 12538
rect 14716 12486 14728 12538
rect 14780 12486 21436 12538
rect 1104 12464 21436 12486
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 9088 12260 10701 12288
rect 9088 12248 9094 12260
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 13814 12288 13820 12300
rect 11011 12260 13820 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 12526 12220 12532 12232
rect 8812 12192 12532 12220
rect 8812 12180 8818 12192
rect 12526 12180 12532 12192
rect 12584 12220 12590 12232
rect 16666 12220 16672 12232
rect 12584 12192 16672 12220
rect 12584 12180 12590 12192
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 16758 12152 16764 12164
rect 11756 12124 16764 12152
rect 11756 12112 11762 12124
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 10870 12084 10876 12096
rect 2832 12056 10876 12084
rect 2832 12044 2838 12056
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 12066 12084 12072 12096
rect 12027 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 1104 11994 21436 12016
rect 1104 11942 4370 11994
rect 4422 11942 4434 11994
rect 4486 11942 4498 11994
rect 4550 11942 4562 11994
rect 4614 11942 11148 11994
rect 11200 11942 11212 11994
rect 11264 11942 11276 11994
rect 11328 11942 11340 11994
rect 11392 11942 17925 11994
rect 17977 11942 17989 11994
rect 18041 11942 18053 11994
rect 18105 11942 18117 11994
rect 18169 11942 21436 11994
rect 1104 11920 21436 11942
rect 3513 11883 3571 11889
rect 3513 11849 3525 11883
rect 3559 11880 3571 11883
rect 9122 11880 9128 11892
rect 3559 11852 9128 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 9122 11840 9128 11852
rect 9180 11880 9186 11892
rect 11882 11880 11888 11892
rect 9180 11852 11888 11880
rect 9180 11840 9186 11852
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 12710 11880 12716 11892
rect 12308 11852 12716 11880
rect 12308 11840 12314 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 13044 11852 16221 11880
rect 13044 11840 13050 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 18322 11812 18328 11824
rect 5040 11784 18328 11812
rect 5040 11772 5046 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 12250 11744 12256 11756
rect 9548 11716 12256 11744
rect 9548 11704 9554 11716
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3620 11648 3801 11676
rect 3142 11568 3148 11620
rect 3200 11608 3206 11620
rect 3620 11608 3648 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 8662 11676 8668 11688
rect 8623 11648 8668 11676
rect 3789 11639 3847 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 10318 11676 10324 11688
rect 9732 11648 10324 11676
rect 9732 11636 9738 11648
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 12710 11676 12716 11688
rect 12667 11648 12716 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 13188 11676 13216 11704
rect 16114 11676 16120 11688
rect 12820 11648 13216 11676
rect 16075 11648 16120 11676
rect 12820 11620 12848 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 3200 11580 3648 11608
rect 3697 11611 3755 11617
rect 3200 11568 3206 11580
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 12342 11608 12348 11620
rect 3743 11580 12348 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 12437 11611 12495 11617
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 12526 11608 12532 11620
rect 12483 11580 12532 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12802 11608 12808 11620
rect 12715 11580 12808 11608
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13170 11608 13176 11620
rect 13131 11580 13176 11608
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 15930 11608 15936 11620
rect 13688 11580 15936 11608
rect 13688 11568 13694 11580
rect 15930 11568 15936 11580
rect 15988 11568 15994 11620
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9582 11540 9588 11552
rect 9088 11512 9588 11540
rect 9088 11500 9094 11512
rect 9582 11500 9588 11512
rect 9640 11540 9646 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9640 11512 9965 11540
rect 9640 11500 9646 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 10376 11512 12725 11540
rect 10376 11500 10382 11512
rect 12713 11509 12725 11512
rect 12759 11540 12771 11543
rect 16574 11540 16580 11552
rect 12759 11512 16580 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 16574 11500 16580 11512
rect 16632 11500 16638 11552
rect 1104 11450 21436 11472
rect 1104 11398 7759 11450
rect 7811 11398 7823 11450
rect 7875 11398 7887 11450
rect 7939 11398 7951 11450
rect 8003 11398 14536 11450
rect 14588 11398 14600 11450
rect 14652 11398 14664 11450
rect 14716 11398 14728 11450
rect 14780 11398 21436 11450
rect 1104 11376 21436 11398
rect 4982 11336 4988 11348
rect 4943 11308 4988 11336
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7650 11336 7656 11348
rect 6963 11308 7656 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9548 11308 10824 11336
rect 9548 11296 9554 11308
rect 4341 11271 4399 11277
rect 4341 11237 4353 11271
rect 4387 11268 4399 11271
rect 6730 11268 6736 11280
rect 4387 11240 6736 11268
rect 4387 11237 4399 11240
rect 4341 11231 4399 11237
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 6822 11228 6828 11280
rect 6880 11228 6886 11280
rect 8754 11268 8760 11280
rect 7576 11240 8760 11268
rect 4571 11203 4629 11209
rect 4571 11169 4583 11203
rect 4617 11200 4629 11203
rect 6840 11200 6868 11228
rect 7576 11209 7604 11240
rect 8754 11228 8760 11240
rect 8812 11268 8818 11280
rect 9398 11268 9404 11280
rect 8812 11240 9404 11268
rect 8812 11228 8818 11240
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 10796 11268 10824 11308
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10928 11308 11069 11336
rect 10928 11296 10934 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 13170 11268 13176 11280
rect 10796 11240 13176 11268
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 4617 11172 6776 11200
rect 6840 11172 6929 11200
rect 4617 11169 4629 11172
rect 4571 11163 4629 11169
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 1820 11104 4721 11132
rect 1820 11092 1826 11104
rect 4709 11101 4721 11104
rect 4755 11132 4767 11135
rect 6748 11132 6776 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 11698 11200 11704 11212
rect 7883 11172 11704 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 8938 11132 8944 11144
rect 4755 11104 6684 11132
rect 6748 11104 8944 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 6656 11064 6684 11104
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 9858 11132 9864 11144
rect 9723 11104 9864 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 9999 11104 18000 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 12066 11064 12072 11076
rect 6656 11036 9720 11064
rect 4506 10999 4564 11005
rect 4506 10965 4518 10999
rect 4552 10996 4564 10999
rect 4706 10996 4712 11008
rect 4552 10968 4712 10996
rect 4552 10965 4564 10968
rect 4506 10959 4564 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8846 10996 8852 11008
rect 8536 10968 8852 10996
rect 8536 10956 8542 10968
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9692 10996 9720 11036
rect 10612 11036 12072 11064
rect 10612 10996 10640 11036
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 9692 10968 10640 10996
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 15194 10996 15200 11008
rect 11572 10968 15200 10996
rect 11572 10956 11578 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 17972 10996 18000 11104
rect 19886 10996 19892 11008
rect 17972 10968 19892 10996
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 1104 10906 21436 10928
rect 1104 10854 4370 10906
rect 4422 10854 4434 10906
rect 4486 10854 4498 10906
rect 4550 10854 4562 10906
rect 4614 10854 11148 10906
rect 11200 10854 11212 10906
rect 11264 10854 11276 10906
rect 11328 10854 11340 10906
rect 11392 10854 17925 10906
rect 17977 10854 17989 10906
rect 18041 10854 18053 10906
rect 18105 10854 18117 10906
rect 18169 10854 21436 10906
rect 1104 10832 21436 10854
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 2648 10764 19840 10792
rect 2648 10752 2654 10764
rect 11514 10724 11520 10736
rect 7116 10696 11520 10724
rect 7116 10597 7144 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 19518 10724 19524 10736
rect 14424 10696 19524 10724
rect 14424 10684 14430 10696
rect 19518 10684 19524 10696
rect 19576 10684 19582 10736
rect 8478 10656 8484 10668
rect 7300 10628 8484 10656
rect 7300 10597 7328 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 9401 10659 9459 10665
rect 8680 10628 9352 10656
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 8680 10588 8708 10628
rect 7699 10560 8708 10588
rect 8941 10591 8999 10597
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9324 10588 9352 10628
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 13906 10656 13912 10668
rect 9447 10628 13912 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 17402 10656 17408 10668
rect 16224 10628 17408 10656
rect 12710 10588 12716 10600
rect 8987 10560 9260 10588
rect 9324 10560 12716 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 8662 10520 8668 10532
rect 8623 10492 8668 10520
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 8849 10523 8907 10529
rect 8849 10520 8861 10523
rect 8812 10492 8861 10520
rect 8812 10480 8818 10492
rect 8849 10489 8861 10492
rect 8895 10489 8907 10523
rect 8849 10483 8907 10489
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10489 9091 10523
rect 9033 10483 9091 10489
rect 2682 10412 2688 10464
rect 2740 10452 2746 10464
rect 9048 10452 9076 10483
rect 9122 10452 9128 10464
rect 2740 10424 9128 10452
rect 2740 10412 2746 10424
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9232 10452 9260 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 16224 10588 16252 10628
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 13219 10560 16252 10588
rect 16301 10591 16359 10597
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 16390 10588 16396 10600
rect 16347 10560 16396 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 16390 10548 16396 10560
rect 16448 10588 16454 10600
rect 17126 10588 17132 10600
rect 16448 10560 17132 10588
rect 16448 10548 16454 10560
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 19610 10588 19616 10600
rect 19571 10560 19616 10588
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 19812 10597 19840 10764
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20073 10795 20131 10801
rect 20073 10792 20085 10795
rect 19944 10764 20085 10792
rect 19944 10752 19950 10764
rect 20073 10761 20085 10764
rect 20119 10761 20131 10795
rect 20073 10755 20131 10761
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10557 19947 10591
rect 19889 10551 19947 10557
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 9364 10492 12296 10520
rect 9364 10480 9370 10492
rect 12268 10464 12296 10492
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 15712 10492 16129 10520
rect 15712 10480 15718 10492
rect 16117 10489 16129 10492
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 16669 10523 16727 10529
rect 16669 10489 16681 10523
rect 16715 10520 16727 10523
rect 18230 10520 18236 10532
rect 16715 10492 18236 10520
rect 16715 10489 16727 10492
rect 16669 10483 16727 10489
rect 18230 10480 18236 10492
rect 18288 10520 18294 10532
rect 18414 10520 18420 10532
rect 18288 10492 18420 10520
rect 18288 10480 18294 10492
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 9674 10452 9680 10464
rect 9232 10424 9680 10452
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 12308 10424 14289 10452
rect 12308 10412 12314 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14277 10415 14335 10421
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 19904 10452 19932 10551
rect 18380 10424 19932 10452
rect 18380 10412 18386 10424
rect 1104 10362 21436 10384
rect 1104 10310 7759 10362
rect 7811 10310 7823 10362
rect 7875 10310 7887 10362
rect 7939 10310 7951 10362
rect 8003 10310 14536 10362
rect 14588 10310 14600 10362
rect 14652 10310 14664 10362
rect 14716 10310 14728 10362
rect 14780 10310 21436 10362
rect 1104 10288 21436 10310
rect 14182 10248 14188 10260
rect 4816 10220 14188 10248
rect 2682 10180 2688 10192
rect 1688 10152 2688 10180
rect 1688 10121 1716 10152
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 4062 10112 4068 10124
rect 1995 10084 4068 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 2409 10047 2467 10053
rect 1452 10016 1900 10044
rect 1452 10004 1458 10016
rect 1762 9976 1768 9988
rect 1723 9948 1768 9976
rect 1762 9936 1768 9948
rect 1820 9936 1826 9988
rect 1872 9976 1900 10016
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 4816 10044 4844 10220
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 15896 10220 17356 10248
rect 15896 10208 15902 10220
rect 10134 10180 10140 10192
rect 10095 10152 10140 10180
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 17328 10189 17356 10220
rect 16945 10183 17003 10189
rect 16945 10180 16957 10183
rect 10428 10152 16957 10180
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 10045 10115 10103 10121
rect 4948 10084 7696 10112
rect 4948 10072 4954 10084
rect 2455 10016 4844 10044
rect 7668 10044 7696 10084
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 10091 10084 10333 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10428 10044 10456 10152
rect 16945 10149 16957 10152
rect 16991 10149 17003 10183
rect 16945 10143 17003 10149
rect 17313 10183 17371 10189
rect 17313 10149 17325 10183
rect 17359 10149 17371 10183
rect 20254 10180 20260 10192
rect 17313 10143 17371 10149
rect 18892 10152 20260 10180
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 14090 10112 14096 10124
rect 10735 10084 14096 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 14976 10084 16773 10112
rect 14976 10072 14982 10084
rect 16761 10081 16773 10084
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 16853 10115 16911 10121
rect 16853 10081 16865 10115
rect 16899 10112 16911 10115
rect 18892 10112 18920 10152
rect 19352 10121 19380 10152
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 16899 10084 18920 10112
rect 18969 10115 19027 10121
rect 16899 10081 16911 10084
rect 16853 10075 16911 10081
rect 18969 10081 18981 10115
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 16574 10044 16580 10056
rect 7668 10016 10456 10044
rect 16535 10016 16580 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 16868 10044 16896 10075
rect 16942 10044 16948 10056
rect 16868 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 18877 9979 18935 9985
rect 18877 9976 18889 9979
rect 1872 9948 18889 9976
rect 18877 9945 18889 9948
rect 18923 9945 18935 9979
rect 18877 9939 18935 9945
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 10042 9908 10048 9920
rect 6788 9880 10048 9908
rect 6788 9868 6794 9880
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 16482 9908 16488 9920
rect 16356 9880 16488 9908
rect 16356 9868 16362 9880
rect 16482 9868 16488 9880
rect 16540 9908 16546 9920
rect 18984 9908 19012 10075
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19576 10016 19625 10044
rect 19576 10004 19582 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 16540 9880 19012 9908
rect 16540 9868 16546 9880
rect 1104 9818 21436 9840
rect 1104 9766 4370 9818
rect 4422 9766 4434 9818
rect 4486 9766 4498 9818
rect 4550 9766 4562 9818
rect 4614 9766 11148 9818
rect 11200 9766 11212 9818
rect 11264 9766 11276 9818
rect 11328 9766 11340 9818
rect 11392 9766 17925 9818
rect 17977 9766 17989 9818
rect 18041 9766 18053 9818
rect 18105 9766 18117 9818
rect 18169 9766 21436 9818
rect 1104 9744 21436 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 9582 9704 9588 9716
rect 4120 9676 9588 9704
rect 4120 9664 4126 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 18230 9704 18236 9716
rect 10100 9676 18236 9704
rect 10100 9664 10106 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4798 9636 4804 9648
rect 4212 9608 4804 9636
rect 4212 9596 4218 9608
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6822 9636 6828 9648
rect 6604 9608 6828 9636
rect 6604 9596 6610 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 9214 9596 9220 9648
rect 9272 9636 9278 9648
rect 9490 9636 9496 9648
rect 9272 9608 9496 9636
rect 9272 9596 9278 9608
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 12894 9636 12900 9648
rect 9916 9608 12900 9636
rect 9916 9596 9922 9608
rect 12894 9596 12900 9608
rect 12952 9636 12958 9648
rect 13722 9636 13728 9648
rect 12952 9608 13728 9636
rect 12952 9596 12958 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 15562 9636 15568 9648
rect 13964 9608 15568 9636
rect 13964 9596 13970 9608
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 20070 9568 20076 9580
rect 3568 9540 20076 9568
rect 3568 9528 3574 9540
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 12526 9500 12532 9512
rect 11940 9472 12532 9500
rect 11940 9460 11946 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14274 9500 14280 9512
rect 13872 9472 14280 9500
rect 13872 9460 13878 9472
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 16632 9472 19993 9500
rect 16632 9460 16638 9472
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 15286 9432 15292 9444
rect 5040 9404 15292 9432
rect 5040 9392 5046 9404
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 7064 9336 8861 9364
rect 7064 9324 7070 9336
rect 8849 9333 8861 9336
rect 8895 9364 8907 9367
rect 9858 9364 9864 9376
rect 8895 9336 9864 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 19610 9364 19616 9376
rect 12584 9336 19616 9364
rect 12584 9324 12590 9336
rect 19610 9324 19616 9336
rect 19668 9364 19674 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19668 9336 20177 9364
rect 19668 9324 19674 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 1104 9274 21436 9296
rect 1104 9222 7759 9274
rect 7811 9222 7823 9274
rect 7875 9222 7887 9274
rect 7939 9222 7951 9274
rect 8003 9222 14536 9274
rect 14588 9222 14600 9274
rect 14652 9222 14664 9274
rect 14716 9222 14728 9274
rect 14780 9222 21436 9274
rect 1104 9200 21436 9222
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5132 9132 11744 9160
rect 5132 9120 5138 9132
rect 3050 9092 3056 9104
rect 3011 9064 3056 9092
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 11716 9092 11744 9132
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 13596 9132 14412 9160
rect 13596 9120 13602 9132
rect 13814 9092 13820 9104
rect 5592 9064 11652 9092
rect 11716 9064 13820 9092
rect 5592 9052 5598 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 7006 9024 7012 9036
rect 1443 8996 7012 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 9640 8996 9781 9024
rect 9640 8984 9646 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 9024 9919 9027
rect 9950 9024 9956 9036
rect 9907 8996 9956 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 9024 11207 9027
rect 11514 9024 11520 9036
rect 11195 8996 11520 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11624 9024 11652 9064
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 13909 9095 13967 9101
rect 13909 9061 13921 9095
rect 13955 9092 13967 9095
rect 14090 9092 14096 9104
rect 13955 9064 14096 9092
rect 13955 9061 13967 9064
rect 13909 9055 13967 9061
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 14384 9101 14412 9132
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9061 14427 9095
rect 14369 9055 14427 9061
rect 13985 9027 14043 9033
rect 13985 9024 13997 9027
rect 11624 8996 13997 9024
rect 13985 8993 13997 8996
rect 14031 9024 14043 9027
rect 14826 9024 14832 9036
rect 14031 8996 14832 9024
rect 14031 8993 14043 8996
rect 13985 8987 14043 8993
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 3970 8956 3976 8968
rect 1912 8928 3976 8956
rect 1912 8916 1918 8928
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 4304 8928 11253 8956
rect 4304 8916 4310 8928
rect 11241 8925 11253 8928
rect 11287 8956 11299 8959
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 11287 8928 13645 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2464 8860 10088 8888
rect 2464 8848 2470 8860
rect 10060 8829 10088 8860
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 16114 8820 16120 8832
rect 15068 8792 16120 8820
rect 15068 8780 15074 8792
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 1104 8730 21436 8752
rect 1104 8678 4370 8730
rect 4422 8678 4434 8730
rect 4486 8678 4498 8730
rect 4550 8678 4562 8730
rect 4614 8678 11148 8730
rect 11200 8678 11212 8730
rect 11264 8678 11276 8730
rect 11328 8678 11340 8730
rect 11392 8678 17925 8730
rect 17977 8678 17989 8730
rect 18041 8678 18053 8730
rect 18105 8678 18117 8730
rect 18169 8678 21436 8730
rect 1104 8656 21436 8678
rect 3602 8616 3608 8628
rect 3563 8588 3608 8616
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 15010 8616 15016 8628
rect 9640 8588 15016 8616
rect 9640 8576 9646 8588
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15470 8616 15476 8628
rect 15160 8588 15476 8616
rect 15160 8576 15166 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 8386 8548 8392 8560
rect 8347 8520 8392 8548
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 19242 8548 19248 8560
rect 11572 8520 19248 8548
rect 11572 8508 11578 8520
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 12894 8480 12900 8492
rect 1728 8452 12900 8480
rect 1728 8440 1734 8452
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3510 8412 3516 8424
rect 2740 8384 3516 8412
rect 2740 8372 2746 8384
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 7006 8412 7012 8424
rect 6967 8384 7012 8412
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 15120 8412 15148 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15804 8452 15945 8480
rect 15804 8440 15810 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 15120 8384 15209 8412
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15344 8384 15393 8412
rect 15344 8372 15350 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 15528 8384 15573 8412
rect 15528 8372 15534 8384
rect 14090 8304 14096 8356
rect 14148 8344 14154 8356
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 14148 8316 15148 8344
rect 14148 8304 14154 8316
rect 15120 8276 15148 8316
rect 15304 8316 15577 8344
rect 15304 8276 15332 8316
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 15565 8307 15623 8313
rect 15120 8248 15332 8276
rect 1104 8186 21436 8208
rect 1104 8134 7759 8186
rect 7811 8134 7823 8186
rect 7875 8134 7887 8186
rect 7939 8134 7951 8186
rect 8003 8134 14536 8186
rect 14588 8134 14600 8186
rect 14652 8134 14664 8186
rect 14716 8134 14728 8186
rect 14780 8134 21436 8186
rect 1104 8112 21436 8134
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 4172 8044 17325 8072
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4172 7945 4200 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 4706 8004 4712 8016
rect 4663 7976 4712 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 11974 8004 11980 8016
rect 11756 7976 11980 8004
rect 11756 7964 11762 7976
rect 11974 7964 11980 7976
rect 12032 8004 12038 8016
rect 12032 7976 17172 8004
rect 12032 7964 12038 7976
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 16850 7936 16856 7948
rect 12860 7908 16856 7936
rect 12860 7896 12866 7908
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 17144 7945 17172 7976
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 7650 7800 7656 7812
rect 2547 7772 7656 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 7650 7760 7656 7772
rect 7708 7800 7714 7812
rect 9398 7800 9404 7812
rect 7708 7772 9404 7800
rect 7708 7760 7714 7772
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 16942 7800 16948 7812
rect 16903 7772 16948 7800
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 5074 7732 5080 7744
rect 3476 7704 5080 7732
rect 3476 7692 3482 7704
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 1104 7642 21436 7664
rect 1104 7590 4370 7642
rect 4422 7590 4434 7642
rect 4486 7590 4498 7642
rect 4550 7590 4562 7642
rect 4614 7590 11148 7642
rect 11200 7590 11212 7642
rect 11264 7590 11276 7642
rect 11328 7590 11340 7642
rect 11392 7590 17925 7642
rect 17977 7590 17989 7642
rect 18041 7590 18053 7642
rect 18105 7590 18117 7642
rect 18169 7590 21436 7642
rect 1104 7568 21436 7590
rect 11514 7528 11520 7540
rect 3804 7500 11520 7528
rect 3160 7364 3648 7392
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 3050 7324 3056 7336
rect 1443 7296 3056 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3160 7333 3188 7364
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7293 3203 7327
rect 3145 7287 3203 7293
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3418 7324 3424 7336
rect 3375 7296 3424 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3528 7188 3556 7287
rect 3620 7256 3648 7364
rect 3804 7333 3832 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 12492 7500 15485 7528
rect 12492 7488 12498 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 13906 7460 13912 7472
rect 4632 7432 13912 7460
rect 4632 7401 4660 7432
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 11790 7392 11796 7404
rect 10183 7364 11796 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 15654 7392 15660 7404
rect 12728 7364 15660 7392
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 4042 7327 4100 7333
rect 4042 7293 4054 7327
rect 4088 7324 4100 7327
rect 4982 7324 4988 7336
rect 4088 7296 4988 7324
rect 4088 7293 4100 7296
rect 4042 7287 4100 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 6604 7296 9781 7324
rect 6604 7284 6610 7296
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 12728 7324 12756 7364
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 9815 7296 12756 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 12952 7296 15393 7324
rect 12952 7284 12958 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 4246 7256 4252 7268
rect 3620 7228 4252 7256
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 9585 7259 9643 7265
rect 9585 7225 9597 7259
rect 9631 7256 9643 7259
rect 12342 7256 12348 7268
rect 9631 7228 12348 7256
rect 9631 7225 9643 7228
rect 9585 7219 9643 7225
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 15194 7256 15200 7268
rect 15155 7228 15200 7256
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 5534 7188 5540 7200
rect 3528 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7188 5598 7200
rect 6638 7188 6644 7200
rect 5592 7160 6644 7188
rect 5592 7148 5598 7160
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 1104 7098 21436 7120
rect 1104 7046 7759 7098
rect 7811 7046 7823 7098
rect 7875 7046 7887 7098
rect 7939 7046 7951 7098
rect 8003 7046 14536 7098
rect 14588 7046 14600 7098
rect 14652 7046 14664 7098
rect 14716 7046 14728 7098
rect 14780 7046 21436 7098
rect 1104 7024 21436 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 6546 6984 6552 6996
rect 1636 6956 6552 6984
rect 1636 6944 1642 6956
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 6822 6916 6828 6928
rect 2823 6888 6828 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 14918 6916 14924 6928
rect 9640 6888 14924 6916
rect 9640 6876 9646 6888
rect 14918 6876 14924 6888
rect 14976 6876 14982 6928
rect 15838 6876 15844 6928
rect 15896 6876 15902 6928
rect 2038 6848 2044 6860
rect 1999 6820 2044 6848
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 1762 6740 1768 6792
rect 1820 6780 1826 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1820 6752 2145 6780
rect 1820 6740 1826 6752
rect 2133 6749 2145 6752
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2332 6712 2360 6811
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 4028 6820 10241 6848
rect 4028 6808 4034 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10410 6848 10416 6860
rect 10367 6820 10416 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 15286 6848 15292 6860
rect 15247 6820 15292 6848
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15436 6851 15494 6857
rect 15436 6817 15448 6851
rect 15482 6848 15494 6851
rect 15856 6848 15884 6876
rect 15482 6820 15884 6848
rect 15482 6817 15494 6820
rect 15436 6811 15494 6817
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 17828 6820 19441 6848
rect 17828 6808 17834 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19613 6851 19671 6857
rect 19613 6817 19625 6851
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 9214 6780 9220 6792
rect 7331 6752 9220 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16390 6780 16396 6792
rect 15896 6752 16396 6780
rect 15896 6740 15902 6752
rect 16390 6740 16396 6752
rect 16448 6780 16454 6792
rect 19628 6780 19656 6811
rect 16448 6752 19656 6780
rect 16448 6740 16454 6752
rect 2332 6684 6776 6712
rect 6748 6644 6776 6684
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 12400 6684 15577 6712
rect 12400 6672 12406 6684
rect 15565 6681 15577 6684
rect 15611 6712 15623 6715
rect 16298 6712 16304 6724
rect 15611 6684 16304 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 6748 6616 8401 6644
rect 8389 6613 8401 6616
rect 8435 6644 8447 6647
rect 11514 6644 11520 6656
rect 8435 6616 11520 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 11514 6604 11520 6616
rect 11572 6644 11578 6656
rect 11698 6644 11704 6656
rect 11572 6616 11704 6644
rect 11572 6604 11578 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 18230 6604 18236 6656
rect 18288 6644 18294 6656
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 18288 6616 19717 6644
rect 18288 6604 18294 6616
rect 19705 6613 19717 6616
rect 19751 6613 19763 6647
rect 19705 6607 19763 6613
rect 1104 6554 21436 6576
rect 1104 6502 4370 6554
rect 4422 6502 4434 6554
rect 4486 6502 4498 6554
rect 4550 6502 4562 6554
rect 4614 6502 11148 6554
rect 11200 6502 11212 6554
rect 11264 6502 11276 6554
rect 11328 6502 11340 6554
rect 11392 6502 17925 6554
rect 17977 6502 17989 6554
rect 18041 6502 18053 6554
rect 18105 6502 18117 6554
rect 18169 6502 21436 6554
rect 1104 6480 21436 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 15838 6440 15844 6452
rect 2096 6412 15844 6440
rect 2096 6400 2102 6412
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 2590 6372 2596 6384
rect 2551 6344 2596 6372
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 15286 6372 15292 6384
rect 6880 6344 15292 6372
rect 6880 6332 6886 6344
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 15746 6304 15752 6316
rect 5316 6276 15752 6304
rect 5316 6264 5322 6276
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 2958 6236 2964 6248
rect 2832 6208 2877 6236
rect 2919 6208 2964 6236
rect 2832 6196 2838 6208
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 17310 6236 17316 6248
rect 3191 6208 17316 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 14090 6168 14096 6180
rect 4212 6140 14096 6168
rect 4212 6128 4218 6140
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 1104 6010 21436 6032
rect 1104 5958 7759 6010
rect 7811 5958 7823 6010
rect 7875 5958 7887 6010
rect 7939 5958 7951 6010
rect 8003 5958 14536 6010
rect 14588 5958 14600 6010
rect 14652 5958 14664 6010
rect 14716 5958 14728 6010
rect 14780 5958 21436 6010
rect 1104 5936 21436 5958
rect 11517 5899 11575 5905
rect 11517 5865 11529 5899
rect 11563 5896 11575 5899
rect 11606 5896 11612 5908
rect 11563 5868 11612 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 2593 5831 2651 5837
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 3326 5828 3332 5840
rect 2639 5800 3332 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 10873 5831 10931 5837
rect 10873 5797 10885 5831
rect 10919 5828 10931 5831
rect 18414 5828 18420 5840
rect 10919 5800 18420 5828
rect 10919 5797 10931 5800
rect 10873 5791 10931 5797
rect 18414 5788 18420 5800
rect 18472 5788 18478 5840
rect 2682 5720 2688 5772
rect 2740 5769 2746 5772
rect 2740 5763 2763 5769
rect 2751 5729 2763 5763
rect 2740 5723 2763 5729
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 4154 5760 4160 5772
rect 3191 5732 4160 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 2740 5720 2746 5723
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 11020 5763 11078 5769
rect 11020 5729 11032 5763
rect 11066 5760 11078 5763
rect 12158 5760 12164 5772
rect 11066 5732 12164 5760
rect 11066 5729 11078 5732
rect 11020 5723 11078 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 11514 5692 11520 5704
rect 11287 5664 11520 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 2409 5627 2467 5633
rect 2409 5593 2421 5627
rect 2455 5624 2467 5627
rect 10134 5624 10140 5636
rect 2455 5596 10140 5624
rect 2455 5593 2467 5596
rect 2409 5587 2467 5593
rect 10134 5584 10140 5596
rect 10192 5584 10198 5636
rect 11149 5627 11207 5633
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 12066 5624 12072 5636
rect 11195 5596 12072 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 1104 5466 21436 5488
rect 1104 5414 4370 5466
rect 4422 5414 4434 5466
rect 4486 5414 4498 5466
rect 4550 5414 4562 5466
rect 4614 5414 11148 5466
rect 11200 5414 11212 5466
rect 11264 5414 11276 5466
rect 11328 5414 11340 5466
rect 11392 5414 17925 5466
rect 17977 5414 17989 5466
rect 18041 5414 18053 5466
rect 18105 5414 18117 5466
rect 18169 5414 21436 5466
rect 1104 5392 21436 5414
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 18322 5352 18328 5364
rect 17276 5324 18328 5352
rect 17276 5312 17282 5324
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 1104 4922 21436 4944
rect 1104 4870 7759 4922
rect 7811 4870 7823 4922
rect 7875 4870 7887 4922
rect 7939 4870 7951 4922
rect 8003 4870 14536 4922
rect 14588 4870 14600 4922
rect 14652 4870 14664 4922
rect 14716 4870 14728 4922
rect 14780 4870 21436 4922
rect 1104 4848 21436 4870
rect 1489 4811 1547 4817
rect 1489 4777 1501 4811
rect 1535 4808 1547 4811
rect 4890 4808 4896 4820
rect 1535 4780 4896 4808
rect 1535 4777 1547 4780
rect 1489 4771 1547 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 16850 4768 16856 4820
rect 16908 4808 16914 4820
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16908 4780 17325 4808
rect 16908 4768 16914 4780
rect 17313 4777 17325 4780
rect 17359 4777 17371 4811
rect 17313 4771 17371 4777
rect 8386 4740 8392 4752
rect 6472 4712 8392 4740
rect 6472 4681 6500 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 1389 4675 1447 4681
rect 1389 4641 1401 4675
rect 1435 4641 1447 4675
rect 1389 4635 1447 4641
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 1412 4604 1440 4635
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 6604 4644 6837 4672
rect 6604 4632 6610 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 7098 4672 7104 4684
rect 7059 4644 7104 4672
rect 6825 4635 6883 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 7616 4644 16221 4672
rect 7616 4632 7622 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 7926 4604 7932 4616
rect 1412 4576 7932 4604
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 13780 4576 15945 4604
rect 13780 4564 13786 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 1104 4378 21436 4400
rect 1104 4326 4370 4378
rect 4422 4326 4434 4378
rect 4486 4326 4498 4378
rect 4550 4326 4562 4378
rect 4614 4326 11148 4378
rect 11200 4326 11212 4378
rect 11264 4326 11276 4378
rect 11328 4326 11340 4378
rect 11392 4326 17925 4378
rect 17977 4326 17989 4378
rect 18041 4326 18053 4378
rect 18105 4326 18117 4378
rect 18169 4326 21436 4378
rect 1104 4304 21436 4326
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7708 4236 7757 4264
rect 7708 4224 7714 4236
rect 7745 4233 7757 4236
rect 7791 4233 7803 4267
rect 7745 4227 7803 4233
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 14366 4196 14372 4208
rect 7984 4168 14372 4196
rect 7984 4156 7990 4168
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 3142 4128 3148 4140
rect 3103 4100 3148 4128
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3878 4128 3884 4140
rect 3839 4100 3884 4128
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 6822 4128 6828 4140
rect 4172 4100 6828 4128
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 4172 4069 4200 4100
rect 6822 4088 6828 4100
rect 6880 4128 6886 4140
rect 8481 4131 8539 4137
rect 6880 4100 8064 4128
rect 6880 4088 6886 4100
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4890 4060 4896 4072
rect 4387 4032 4896 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 7926 4060 7932 4072
rect 7887 4032 7932 4060
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8036 4069 8064 4100
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8570 4128 8576 4140
rect 8527 4100 8576 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 19150 4128 19156 4140
rect 15988 4100 19156 4128
rect 15988 4088 15994 4100
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 12526 4060 12532 4072
rect 8168 4032 11468 4060
rect 12487 4032 12532 4060
rect 8168 4020 8174 4032
rect 11440 3992 11468 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13446 4060 13452 4072
rect 12851 4032 13452 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13265 3995 13323 4001
rect 13265 3992 13277 3995
rect 11440 3964 13277 3992
rect 13265 3961 13277 3964
rect 13311 3961 13323 3995
rect 13265 3955 13323 3961
rect 1104 3834 21436 3856
rect 1104 3782 7759 3834
rect 7811 3782 7823 3834
rect 7875 3782 7887 3834
rect 7939 3782 7951 3834
rect 8003 3782 14536 3834
rect 14588 3782 14600 3834
rect 14652 3782 14664 3834
rect 14716 3782 14728 3834
rect 14780 3782 21436 3834
rect 1104 3760 21436 3782
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 7340 3692 10793 3720
rect 7340 3680 7346 3692
rect 10781 3689 10793 3692
rect 10827 3689 10839 3723
rect 10781 3683 10839 3689
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 1104 3290 21436 3312
rect 1104 3238 4370 3290
rect 4422 3238 4434 3290
rect 4486 3238 4498 3290
rect 4550 3238 4562 3290
rect 4614 3238 11148 3290
rect 11200 3238 11212 3290
rect 11264 3238 11276 3290
rect 11328 3238 11340 3290
rect 11392 3238 17925 3290
rect 17977 3238 17989 3290
rect 18041 3238 18053 3290
rect 18105 3238 18117 3290
rect 18169 3238 21436 3290
rect 1104 3216 21436 3238
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4304 3012 4445 3040
rect 4304 3000 4310 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 4433 3003 4491 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 4212 2944 4721 2972
rect 4212 2932 4218 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 16172 2944 20085 2972
rect 16172 2932 16178 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 4801 2907 4859 2913
rect 4801 2873 4813 2907
rect 4847 2904 4859 2907
rect 15102 2904 15108 2916
rect 4847 2876 15108 2904
rect 4847 2873 4859 2876
rect 4801 2867 4859 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 4617 2839 4675 2845
rect 4617 2836 4629 2839
rect 624 2808 4629 2836
rect 624 2796 630 2808
rect 4617 2805 4629 2808
rect 4663 2836 4675 2839
rect 5074 2836 5080 2848
rect 4663 2808 5080 2836
rect 4663 2805 4675 2808
rect 4617 2799 4675 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8662 2836 8668 2848
rect 8352 2808 8668 2836
rect 8352 2796 8358 2808
rect 8662 2796 8668 2808
rect 8720 2836 8726 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 8720 2808 20269 2836
rect 8720 2796 8726 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20257 2799 20315 2805
rect 1104 2746 21436 2768
rect 1104 2694 7759 2746
rect 7811 2694 7823 2746
rect 7875 2694 7887 2746
rect 7939 2694 7951 2746
rect 8003 2694 14536 2746
rect 14588 2694 14600 2746
rect 14652 2694 14664 2746
rect 14716 2694 14728 2746
rect 14780 2694 21436 2746
rect 1104 2672 21436 2694
rect 7024 2604 10640 2632
rect 7024 2564 7052 2604
rect 6932 2536 7052 2564
rect 6932 2505 6960 2536
rect 7650 2524 7656 2576
rect 7708 2564 7714 2576
rect 7708 2536 8432 2564
rect 7708 2524 7714 2536
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 8294 2496 8300 2508
rect 7055 2468 8300 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8404 2496 8432 2536
rect 8938 2524 8944 2576
rect 8996 2564 9002 2576
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 8996 2536 10517 2564
rect 8996 2524 9002 2536
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10612 2564 10640 2604
rect 16942 2564 16948 2576
rect 10612 2536 16948 2564
rect 10505 2527 10563 2533
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 8404 2468 11069 2496
rect 11057 2465 11069 2468
rect 11103 2465 11115 2499
rect 11057 2459 11115 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 12250 2496 12256 2508
rect 11563 2468 12256 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 11348 2428 11376 2459
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 7515 2400 11376 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 1104 2202 21436 2224
rect 1104 2150 4370 2202
rect 4422 2150 4434 2202
rect 4486 2150 4498 2202
rect 4550 2150 4562 2202
rect 4614 2150 11148 2202
rect 11200 2150 11212 2202
rect 11264 2150 11276 2202
rect 11328 2150 11340 2202
rect 11392 2150 17925 2202
rect 17977 2150 17989 2202
rect 18041 2150 18053 2202
rect 18105 2150 18117 2202
rect 18169 2150 21436 2202
rect 1104 2128 21436 2150
<< via1 >>
rect 7759 22278 7811 22330
rect 7823 22278 7875 22330
rect 7887 22278 7939 22330
rect 7951 22278 8003 22330
rect 14536 22278 14588 22330
rect 14600 22278 14652 22330
rect 14664 22278 14716 22330
rect 14728 22278 14780 22330
rect 8576 22108 8628 22160
rect 15292 22040 15344 22092
rect 7380 21904 7432 21956
rect 19708 21904 19760 21956
rect 13452 21836 13504 21888
rect 4370 21734 4422 21786
rect 4434 21734 4486 21786
rect 4498 21734 4550 21786
rect 4562 21734 4614 21786
rect 11148 21734 11200 21786
rect 11212 21734 11264 21786
rect 11276 21734 11328 21786
rect 11340 21734 11392 21786
rect 17925 21734 17977 21786
rect 17989 21734 18041 21786
rect 18053 21734 18105 21786
rect 18117 21734 18169 21786
rect 12072 21564 12124 21616
rect 18972 21564 19024 21616
rect 11980 21496 12032 21548
rect 13176 21428 13228 21480
rect 16948 21428 17000 21480
rect 19708 21471 19760 21480
rect 19708 21437 19717 21471
rect 19717 21437 19751 21471
rect 19751 21437 19760 21471
rect 19708 21428 19760 21437
rect 19892 21471 19944 21480
rect 19892 21437 19901 21471
rect 19901 21437 19935 21471
rect 19935 21437 19944 21471
rect 19892 21428 19944 21437
rect 9220 21403 9272 21412
rect 9220 21369 9229 21403
rect 9229 21369 9263 21403
rect 9263 21369 9272 21403
rect 9220 21360 9272 21369
rect 16304 21360 16356 21412
rect 16580 21292 16632 21344
rect 7759 21190 7811 21242
rect 7823 21190 7875 21242
rect 7887 21190 7939 21242
rect 7951 21190 8003 21242
rect 14536 21190 14588 21242
rect 14600 21190 14652 21242
rect 14664 21190 14716 21242
rect 14728 21190 14780 21242
rect 17592 21088 17644 21140
rect 19892 21088 19944 21140
rect 16764 21020 16816 21072
rect 20260 21020 20312 21072
rect 6368 20952 6420 21004
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 16396 20952 16448 21004
rect 10692 20884 10744 20936
rect 16672 20884 16724 20936
rect 8300 20816 8352 20868
rect 17408 20816 17460 20868
rect 4370 20646 4422 20698
rect 4434 20646 4486 20698
rect 4498 20646 4550 20698
rect 4562 20646 4614 20698
rect 11148 20646 11200 20698
rect 11212 20646 11264 20698
rect 11276 20646 11328 20698
rect 11340 20646 11392 20698
rect 17925 20646 17977 20698
rect 17989 20646 18041 20698
rect 18053 20646 18105 20698
rect 18117 20646 18169 20698
rect 9588 20544 9640 20596
rect 12164 20544 12216 20596
rect 12716 20544 12768 20596
rect 12716 20408 12768 20460
rect 14832 20340 14884 20392
rect 17500 20340 17552 20392
rect 8392 20272 8444 20324
rect 15844 20272 15896 20324
rect 15108 20204 15160 20256
rect 17040 20204 17092 20256
rect 19340 20204 19392 20256
rect 7759 20102 7811 20154
rect 7823 20102 7875 20154
rect 7887 20102 7939 20154
rect 7951 20102 8003 20154
rect 14536 20102 14588 20154
rect 14600 20102 14652 20154
rect 14664 20102 14716 20154
rect 14728 20102 14780 20154
rect 10140 20000 10192 20052
rect 2964 19932 3016 19984
rect 8852 19932 8904 19984
rect 21916 19932 21968 19984
rect 11520 19864 11572 19916
rect 16396 19907 16448 19916
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 16672 19864 16724 19916
rect 11796 19796 11848 19848
rect 17592 19796 17644 19848
rect 15016 19660 15068 19712
rect 4370 19558 4422 19610
rect 4434 19558 4486 19610
rect 4498 19558 4550 19610
rect 4562 19558 4614 19610
rect 11148 19558 11200 19610
rect 11212 19558 11264 19610
rect 11276 19558 11328 19610
rect 11340 19558 11392 19610
rect 17925 19558 17977 19610
rect 17989 19558 18041 19610
rect 18053 19558 18105 19610
rect 18117 19558 18169 19610
rect 3332 19320 3384 19372
rect 8668 19320 8720 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 7380 19116 7432 19168
rect 8116 19252 8168 19304
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 13636 19295 13688 19304
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 16488 19184 16540 19236
rect 8484 19116 8536 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 7759 19014 7811 19066
rect 7823 19014 7875 19066
rect 7887 19014 7939 19066
rect 7951 19014 8003 19066
rect 14536 19014 14588 19066
rect 14600 19014 14652 19066
rect 14664 19014 14716 19066
rect 14728 19014 14780 19066
rect 1952 18912 2004 18964
rect 17316 18912 17368 18964
rect 17224 18844 17276 18896
rect 17592 18844 17644 18896
rect 13360 18776 13412 18828
rect 16856 18708 16908 18760
rect 4370 18470 4422 18522
rect 4434 18470 4486 18522
rect 4498 18470 4550 18522
rect 4562 18470 4614 18522
rect 11148 18470 11200 18522
rect 11212 18470 11264 18522
rect 11276 18470 11328 18522
rect 11340 18470 11392 18522
rect 17925 18470 17977 18522
rect 17989 18470 18041 18522
rect 18053 18470 18105 18522
rect 18117 18470 18169 18522
rect 11704 18232 11756 18284
rect 3608 18096 3660 18148
rect 13268 18164 13320 18216
rect 18972 18164 19024 18216
rect 7564 18139 7616 18148
rect 6920 18028 6972 18080
rect 7564 18105 7573 18139
rect 7573 18105 7607 18139
rect 7607 18105 7616 18139
rect 7564 18096 7616 18105
rect 20260 18071 20312 18080
rect 20260 18037 20269 18071
rect 20269 18037 20303 18071
rect 20303 18037 20312 18071
rect 20260 18028 20312 18037
rect 7759 17926 7811 17978
rect 7823 17926 7875 17978
rect 7887 17926 7939 17978
rect 7951 17926 8003 17978
rect 14536 17926 14588 17978
rect 14600 17926 14652 17978
rect 14664 17926 14716 17978
rect 14728 17926 14780 17978
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 12164 17756 12216 17808
rect 14372 17756 14424 17808
rect 10416 17688 10468 17740
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 11612 17620 11664 17672
rect 2688 17552 2740 17604
rect 15660 17552 15712 17604
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 4370 17382 4422 17434
rect 4434 17382 4486 17434
rect 4498 17382 4550 17434
rect 4562 17382 4614 17434
rect 11148 17382 11200 17434
rect 11212 17382 11264 17434
rect 11276 17382 11328 17434
rect 11340 17382 11392 17434
rect 17925 17382 17977 17434
rect 17989 17382 18041 17434
rect 18053 17382 18105 17434
rect 18117 17382 18169 17434
rect 17040 17280 17092 17332
rect 5356 17144 5408 17196
rect 13084 17144 13136 17196
rect 5264 17076 5316 17128
rect 6736 17076 6788 17128
rect 3792 17008 3844 17060
rect 15292 17008 15344 17060
rect 9496 16940 9548 16992
rect 16396 16940 16448 16992
rect 7759 16838 7811 16890
rect 7823 16838 7875 16890
rect 7887 16838 7939 16890
rect 7951 16838 8003 16890
rect 14536 16838 14588 16890
rect 14600 16838 14652 16890
rect 14664 16838 14716 16890
rect 14728 16838 14780 16890
rect 14004 16736 14056 16788
rect 11704 16668 11756 16720
rect 2964 16600 3016 16652
rect 12992 16643 13044 16652
rect 12992 16609 13001 16643
rect 13001 16609 13035 16643
rect 13035 16609 13044 16643
rect 12992 16600 13044 16609
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 16580 16668 16632 16720
rect 16856 16711 16908 16720
rect 16856 16677 16865 16711
rect 16865 16677 16899 16711
rect 16899 16677 16908 16711
rect 16856 16668 16908 16677
rect 16580 16532 16632 16584
rect 16764 16532 16816 16584
rect 4370 16294 4422 16346
rect 4434 16294 4486 16346
rect 4498 16294 4550 16346
rect 4562 16294 4614 16346
rect 11148 16294 11200 16346
rect 11212 16294 11264 16346
rect 11276 16294 11328 16346
rect 11340 16294 11392 16346
rect 17925 16294 17977 16346
rect 17989 16294 18041 16346
rect 18053 16294 18105 16346
rect 18117 16294 18169 16346
rect 6736 16192 6788 16244
rect 14280 16235 14332 16244
rect 14280 16201 14289 16235
rect 14289 16201 14323 16235
rect 14323 16201 14332 16235
rect 14280 16192 14332 16201
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 2412 15920 2464 15972
rect 2688 15920 2740 15972
rect 7104 15988 7156 16040
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 7656 16031 7708 16040
rect 7656 15997 7665 16031
rect 7665 15997 7699 16031
rect 7699 15997 7708 16031
rect 7656 15988 7708 15997
rect 8300 15920 8352 15972
rect 6736 15852 6788 15904
rect 9956 15852 10008 15904
rect 14188 15988 14240 16040
rect 7759 15750 7811 15802
rect 7823 15750 7875 15802
rect 7887 15750 7939 15802
rect 7951 15750 8003 15802
rect 14536 15750 14588 15802
rect 14600 15750 14652 15802
rect 14664 15750 14716 15802
rect 14728 15750 14780 15802
rect 2872 15580 2924 15632
rect 13728 15580 13780 15632
rect 5080 15512 5132 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 15200 15308 15252 15360
rect 4370 15206 4422 15258
rect 4434 15206 4486 15258
rect 4498 15206 4550 15258
rect 4562 15206 4614 15258
rect 11148 15206 11200 15258
rect 11212 15206 11264 15258
rect 11276 15206 11328 15258
rect 11340 15206 11392 15258
rect 17925 15206 17977 15258
rect 17989 15206 18041 15258
rect 18053 15206 18105 15258
rect 18117 15206 18169 15258
rect 11520 14968 11572 15020
rect 13176 14968 13228 15020
rect 3516 14943 3568 14952
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 4252 14900 4304 14952
rect 14280 14968 14332 15020
rect 13912 14900 13964 14952
rect 14096 14832 14148 14884
rect 15844 14832 15896 14884
rect 12440 14764 12492 14816
rect 13820 14764 13872 14816
rect 7759 14662 7811 14714
rect 7823 14662 7875 14714
rect 7887 14662 7939 14714
rect 7951 14662 8003 14714
rect 14536 14662 14588 14714
rect 14600 14662 14652 14714
rect 14664 14662 14716 14714
rect 14728 14662 14780 14714
rect 3240 14560 3292 14612
rect 3516 14560 3568 14612
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 9036 14560 9088 14612
rect 9588 14424 9640 14476
rect 10048 14560 10100 14612
rect 19340 14560 19392 14612
rect 13084 14492 13136 14544
rect 17040 14424 17092 14476
rect 18236 14424 18288 14476
rect 5172 14356 5224 14408
rect 4068 14220 4120 14272
rect 13268 14356 13320 14408
rect 17316 14356 17368 14408
rect 17776 14356 17828 14408
rect 9680 14220 9732 14272
rect 4370 14118 4422 14170
rect 4434 14118 4486 14170
rect 4498 14118 4550 14170
rect 4562 14118 4614 14170
rect 11148 14118 11200 14170
rect 11212 14118 11264 14170
rect 11276 14118 11328 14170
rect 11340 14118 11392 14170
rect 17925 14118 17977 14170
rect 17989 14118 18041 14170
rect 18053 14118 18105 14170
rect 18117 14118 18169 14170
rect 7759 13574 7811 13626
rect 7823 13574 7875 13626
rect 7887 13574 7939 13626
rect 7951 13574 8003 13626
rect 14536 13574 14588 13626
rect 14600 13574 14652 13626
rect 14664 13574 14716 13626
rect 14728 13574 14780 13626
rect 17316 13472 17368 13524
rect 17500 13515 17552 13524
rect 17500 13481 17509 13515
rect 17509 13481 17543 13515
rect 17543 13481 17552 13515
rect 17500 13472 17552 13481
rect 16764 13404 16816 13456
rect 16948 13404 17000 13456
rect 6920 13336 6972 13388
rect 3884 13268 3936 13320
rect 13636 13268 13688 13320
rect 16488 13336 16540 13388
rect 17132 13336 17184 13388
rect 3056 13200 3108 13252
rect 13452 13132 13504 13184
rect 15384 13132 15436 13184
rect 4370 13030 4422 13082
rect 4434 13030 4486 13082
rect 4498 13030 4550 13082
rect 4562 13030 4614 13082
rect 11148 13030 11200 13082
rect 11212 13030 11264 13082
rect 11276 13030 11328 13082
rect 11340 13030 11392 13082
rect 17925 13030 17977 13082
rect 17989 13030 18041 13082
rect 18053 13030 18105 13082
rect 18117 13030 18169 13082
rect 3424 12928 3476 12980
rect 6920 12928 6972 12980
rect 13636 12928 13688 12980
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 13452 12860 13504 12912
rect 14096 12860 14148 12912
rect 14924 12860 14976 12912
rect 11796 12724 11848 12776
rect 14280 12724 14332 12776
rect 19248 12792 19300 12844
rect 15108 12724 15160 12776
rect 14372 12699 14424 12708
rect 14372 12665 14381 12699
rect 14381 12665 14415 12699
rect 14415 12665 14424 12699
rect 14372 12656 14424 12665
rect 15016 12656 15068 12708
rect 9128 12588 9180 12640
rect 11704 12588 11756 12640
rect 14004 12588 14056 12640
rect 14280 12588 14332 12640
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 7759 12486 7811 12538
rect 7823 12486 7875 12538
rect 7887 12486 7939 12538
rect 7951 12486 8003 12538
rect 14536 12486 14588 12538
rect 14600 12486 14652 12538
rect 14664 12486 14716 12538
rect 14728 12486 14780 12538
rect 9036 12248 9088 12300
rect 13820 12248 13872 12300
rect 8760 12180 8812 12232
rect 12532 12180 12584 12232
rect 16672 12180 16724 12232
rect 11704 12112 11756 12164
rect 16764 12112 16816 12164
rect 2780 12044 2832 12096
rect 10876 12044 10928 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 4370 11942 4422 11994
rect 4434 11942 4486 11994
rect 4498 11942 4550 11994
rect 4562 11942 4614 11994
rect 11148 11942 11200 11994
rect 11212 11942 11264 11994
rect 11276 11942 11328 11994
rect 11340 11942 11392 11994
rect 17925 11942 17977 11994
rect 17989 11942 18041 11994
rect 18053 11942 18105 11994
rect 18117 11942 18169 11994
rect 9128 11840 9180 11892
rect 11888 11840 11940 11892
rect 12256 11840 12308 11892
rect 12716 11840 12768 11892
rect 12992 11840 13044 11892
rect 4988 11772 5040 11824
rect 18328 11772 18380 11824
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 9496 11704 9548 11756
rect 12256 11704 12308 11756
rect 13176 11704 13228 11756
rect 3148 11568 3200 11620
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9680 11636 9732 11688
rect 10324 11636 10376 11688
rect 12716 11636 12768 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 12348 11568 12400 11620
rect 12532 11568 12584 11620
rect 12808 11611 12860 11620
rect 12808 11577 12817 11611
rect 12817 11577 12851 11611
rect 12851 11577 12860 11611
rect 12808 11568 12860 11577
rect 13176 11611 13228 11620
rect 13176 11577 13185 11611
rect 13185 11577 13219 11611
rect 13219 11577 13228 11611
rect 13176 11568 13228 11577
rect 13636 11568 13688 11620
rect 15936 11611 15988 11620
rect 15936 11577 15945 11611
rect 15945 11577 15979 11611
rect 15979 11577 15988 11611
rect 15936 11568 15988 11577
rect 9036 11500 9088 11552
rect 9588 11500 9640 11552
rect 10324 11500 10376 11552
rect 16580 11500 16632 11552
rect 7759 11398 7811 11450
rect 7823 11398 7875 11450
rect 7887 11398 7939 11450
rect 7951 11398 8003 11450
rect 14536 11398 14588 11450
rect 14600 11398 14652 11450
rect 14664 11398 14716 11450
rect 14728 11398 14780 11450
rect 4988 11339 5040 11348
rect 4988 11305 4997 11339
rect 4997 11305 5031 11339
rect 5031 11305 5040 11339
rect 4988 11296 5040 11305
rect 7656 11296 7708 11348
rect 9496 11296 9548 11348
rect 6736 11228 6788 11280
rect 6828 11228 6880 11280
rect 8760 11228 8812 11280
rect 9404 11228 9456 11280
rect 10876 11296 10928 11348
rect 13176 11228 13228 11280
rect 1768 11092 1820 11144
rect 11704 11160 11756 11212
rect 8944 11092 8996 11144
rect 9864 11092 9916 11144
rect 4712 10956 4764 11008
rect 8484 10956 8536 11008
rect 8852 10956 8904 11008
rect 12072 11024 12124 11076
rect 11520 10956 11572 11008
rect 15200 10956 15252 11008
rect 19892 10956 19944 11008
rect 4370 10854 4422 10906
rect 4434 10854 4486 10906
rect 4498 10854 4550 10906
rect 4562 10854 4614 10906
rect 11148 10854 11200 10906
rect 11212 10854 11264 10906
rect 11276 10854 11328 10906
rect 11340 10854 11392 10906
rect 17925 10854 17977 10906
rect 17989 10854 18041 10906
rect 18053 10854 18105 10906
rect 18117 10854 18169 10906
rect 2596 10752 2648 10804
rect 11520 10684 11572 10736
rect 14372 10684 14424 10736
rect 19524 10684 19576 10736
rect 8484 10616 8536 10668
rect 13912 10616 13964 10668
rect 8668 10523 8720 10532
rect 8668 10489 8677 10523
rect 8677 10489 8711 10523
rect 8711 10489 8720 10523
rect 8668 10480 8720 10489
rect 8760 10480 8812 10532
rect 2688 10412 2740 10464
rect 9128 10412 9180 10464
rect 12716 10548 12768 10600
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 17408 10616 17460 10668
rect 16396 10548 16448 10600
rect 17132 10548 17184 10600
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 19892 10752 19944 10804
rect 9312 10480 9364 10532
rect 15660 10480 15712 10532
rect 18236 10480 18288 10532
rect 18420 10480 18472 10532
rect 9680 10412 9732 10464
rect 12256 10412 12308 10464
rect 18328 10412 18380 10464
rect 7759 10310 7811 10362
rect 7823 10310 7875 10362
rect 7887 10310 7939 10362
rect 7951 10310 8003 10362
rect 14536 10310 14588 10362
rect 14600 10310 14652 10362
rect 14664 10310 14716 10362
rect 14728 10310 14780 10362
rect 2688 10140 2740 10192
rect 4068 10072 4120 10124
rect 1400 10004 1452 10056
rect 1768 9979 1820 9988
rect 1768 9945 1777 9979
rect 1777 9945 1811 9979
rect 1811 9945 1820 9979
rect 1768 9936 1820 9945
rect 14188 10208 14240 10260
rect 15844 10208 15896 10260
rect 10140 10183 10192 10192
rect 10140 10149 10149 10183
rect 10149 10149 10183 10183
rect 10183 10149 10192 10183
rect 10140 10140 10192 10149
rect 4896 10072 4948 10124
rect 14096 10072 14148 10124
rect 14924 10072 14976 10124
rect 20260 10140 20312 10192
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 16948 10004 17000 10056
rect 6736 9868 6788 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 16304 9868 16356 9920
rect 16488 9868 16540 9920
rect 19524 10004 19576 10056
rect 4370 9766 4422 9818
rect 4434 9766 4486 9818
rect 4498 9766 4550 9818
rect 4562 9766 4614 9818
rect 11148 9766 11200 9818
rect 11212 9766 11264 9818
rect 11276 9766 11328 9818
rect 11340 9766 11392 9818
rect 17925 9766 17977 9818
rect 17989 9766 18041 9818
rect 18053 9766 18105 9818
rect 18117 9766 18169 9818
rect 4068 9664 4120 9716
rect 9588 9664 9640 9716
rect 10048 9664 10100 9716
rect 18236 9664 18288 9716
rect 4160 9596 4212 9648
rect 4804 9596 4856 9648
rect 6552 9596 6604 9648
rect 6828 9596 6880 9648
rect 9220 9596 9272 9648
rect 9496 9596 9548 9648
rect 9864 9596 9916 9648
rect 12900 9596 12952 9648
rect 13728 9596 13780 9648
rect 13912 9596 13964 9648
rect 15568 9596 15620 9648
rect 3516 9528 3568 9580
rect 20076 9528 20128 9580
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 11888 9460 11940 9512
rect 12532 9460 12584 9512
rect 13820 9460 13872 9512
rect 14280 9460 14332 9512
rect 16580 9460 16632 9512
rect 4988 9392 5040 9444
rect 15292 9392 15344 9444
rect 7012 9324 7064 9376
rect 9864 9324 9916 9376
rect 12532 9324 12584 9376
rect 19616 9324 19668 9376
rect 7759 9222 7811 9274
rect 7823 9222 7875 9274
rect 7887 9222 7939 9274
rect 7951 9222 8003 9274
rect 14536 9222 14588 9274
rect 14600 9222 14652 9274
rect 14664 9222 14716 9274
rect 14728 9222 14780 9274
rect 5080 9120 5132 9172
rect 3056 9095 3108 9104
rect 3056 9061 3065 9095
rect 3065 9061 3099 9095
rect 3099 9061 3108 9095
rect 3056 9052 3108 9061
rect 5540 9052 5592 9104
rect 13544 9120 13596 9172
rect 13820 9095 13872 9104
rect 7012 8984 7064 9036
rect 9588 8984 9640 9036
rect 9956 8984 10008 9036
rect 11520 8984 11572 9036
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 14096 9052 14148 9104
rect 14832 8984 14884 9036
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 1860 8916 1912 8968
rect 3976 8916 4028 8968
rect 4252 8916 4304 8968
rect 2412 8848 2464 8900
rect 15016 8780 15068 8832
rect 16120 8780 16172 8832
rect 4370 8678 4422 8730
rect 4434 8678 4486 8730
rect 4498 8678 4550 8730
rect 4562 8678 4614 8730
rect 11148 8678 11200 8730
rect 11212 8678 11264 8730
rect 11276 8678 11328 8730
rect 11340 8678 11392 8730
rect 17925 8678 17977 8730
rect 17989 8678 18041 8730
rect 18053 8678 18105 8730
rect 18117 8678 18169 8730
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 9588 8576 9640 8628
rect 15016 8576 15068 8628
rect 15108 8576 15160 8628
rect 15476 8576 15528 8628
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 11520 8508 11572 8560
rect 1676 8440 1728 8492
rect 12900 8440 12952 8492
rect 2688 8372 2740 8424
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 19248 8508 19300 8560
rect 15752 8440 15804 8492
rect 15292 8372 15344 8424
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 14096 8304 14148 8356
rect 7759 8134 7811 8186
rect 7823 8134 7875 8186
rect 7887 8134 7939 8186
rect 7951 8134 8003 8186
rect 14536 8134 14588 8186
rect 14600 8134 14652 8186
rect 14664 8134 14716 8186
rect 14728 8134 14780 8186
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4712 7964 4764 8016
rect 11704 7964 11756 8016
rect 11980 7964 12032 8016
rect 12808 7896 12860 7948
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 7656 7760 7708 7812
rect 9404 7760 9456 7812
rect 16948 7803 17000 7812
rect 16948 7769 16957 7803
rect 16957 7769 16991 7803
rect 16991 7769 17000 7803
rect 16948 7760 17000 7769
rect 3424 7692 3476 7744
rect 5080 7692 5132 7744
rect 4370 7590 4422 7642
rect 4434 7590 4486 7642
rect 4498 7590 4550 7642
rect 4562 7590 4614 7642
rect 11148 7590 11200 7642
rect 11212 7590 11264 7642
rect 11276 7590 11328 7642
rect 11340 7590 11392 7642
rect 17925 7590 17977 7642
rect 17989 7590 18041 7642
rect 18053 7590 18105 7642
rect 18117 7590 18169 7642
rect 3056 7284 3108 7336
rect 3424 7284 3476 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 11520 7488 11572 7540
rect 12440 7488 12492 7540
rect 13912 7420 13964 7472
rect 11796 7352 11848 7404
rect 4988 7284 5040 7336
rect 6552 7284 6604 7336
rect 15660 7352 15712 7404
rect 12900 7284 12952 7336
rect 4252 7216 4304 7268
rect 12348 7216 12400 7268
rect 15200 7259 15252 7268
rect 15200 7225 15209 7259
rect 15209 7225 15243 7259
rect 15243 7225 15252 7259
rect 15200 7216 15252 7225
rect 5540 7148 5592 7200
rect 6644 7148 6696 7200
rect 7759 7046 7811 7098
rect 7823 7046 7875 7098
rect 7887 7046 7939 7098
rect 7951 7046 8003 7098
rect 14536 7046 14588 7098
rect 14600 7046 14652 7098
rect 14664 7046 14716 7098
rect 14728 7046 14780 7098
rect 1584 6944 1636 6996
rect 6552 6944 6604 6996
rect 6828 6876 6880 6928
rect 9588 6876 9640 6928
rect 14924 6876 14976 6928
rect 15844 6876 15896 6928
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 1768 6740 1820 6792
rect 3976 6808 4028 6860
rect 10416 6808 10468 6860
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 17776 6808 17828 6860
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 9220 6740 9272 6792
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 15844 6740 15896 6792
rect 16396 6740 16448 6792
rect 12348 6672 12400 6724
rect 16304 6672 16356 6724
rect 11520 6604 11572 6656
rect 11704 6604 11756 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 18236 6604 18288 6656
rect 4370 6502 4422 6554
rect 4434 6502 4486 6554
rect 4498 6502 4550 6554
rect 4562 6502 4614 6554
rect 11148 6502 11200 6554
rect 11212 6502 11264 6554
rect 11276 6502 11328 6554
rect 11340 6502 11392 6554
rect 17925 6502 17977 6554
rect 17989 6502 18041 6554
rect 18053 6502 18105 6554
rect 18117 6502 18169 6554
rect 2044 6400 2096 6452
rect 15844 6400 15896 6452
rect 2596 6375 2648 6384
rect 2596 6341 2605 6375
rect 2605 6341 2639 6375
rect 2639 6341 2648 6375
rect 2596 6332 2648 6341
rect 6828 6332 6880 6384
rect 15292 6332 15344 6384
rect 5264 6264 5316 6316
rect 15752 6264 15804 6316
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2964 6239 3016 6248
rect 2780 6196 2832 6205
rect 2964 6205 2973 6239
rect 2973 6205 3007 6239
rect 3007 6205 3016 6239
rect 2964 6196 3016 6205
rect 17316 6196 17368 6248
rect 4160 6128 4212 6180
rect 14096 6128 14148 6180
rect 7759 5958 7811 6010
rect 7823 5958 7875 6010
rect 7887 5958 7939 6010
rect 7951 5958 8003 6010
rect 14536 5958 14588 6010
rect 14600 5958 14652 6010
rect 14664 5958 14716 6010
rect 14728 5958 14780 6010
rect 11612 5856 11664 5908
rect 3332 5788 3384 5840
rect 18420 5788 18472 5840
rect 2688 5763 2740 5772
rect 2688 5729 2717 5763
rect 2717 5729 2740 5763
rect 2688 5720 2740 5729
rect 4160 5720 4212 5772
rect 12164 5720 12216 5772
rect 11520 5652 11572 5704
rect 10140 5584 10192 5636
rect 12072 5584 12124 5636
rect 4370 5414 4422 5466
rect 4434 5414 4486 5466
rect 4498 5414 4550 5466
rect 4562 5414 4614 5466
rect 11148 5414 11200 5466
rect 11212 5414 11264 5466
rect 11276 5414 11328 5466
rect 11340 5414 11392 5466
rect 17925 5414 17977 5466
rect 17989 5414 18041 5466
rect 18053 5414 18105 5466
rect 18117 5414 18169 5466
rect 17224 5312 17276 5364
rect 18328 5312 18380 5364
rect 7759 4870 7811 4922
rect 7823 4870 7875 4922
rect 7887 4870 7939 4922
rect 7951 4870 8003 4922
rect 14536 4870 14588 4922
rect 14600 4870 14652 4922
rect 14664 4870 14716 4922
rect 14728 4870 14780 4922
rect 4896 4768 4948 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 16856 4768 16908 4820
rect 8392 4700 8444 4752
rect 6552 4632 6604 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7564 4632 7616 4684
rect 7932 4564 7984 4616
rect 13728 4564 13780 4616
rect 4370 4326 4422 4378
rect 4434 4326 4486 4378
rect 4498 4326 4550 4378
rect 4562 4326 4614 4378
rect 11148 4326 11200 4378
rect 11212 4326 11264 4378
rect 11276 4326 11328 4378
rect 11340 4326 11392 4378
rect 17925 4326 17977 4378
rect 17989 4326 18041 4378
rect 18053 4326 18105 4378
rect 18117 4326 18169 4378
rect 7656 4224 7708 4276
rect 7932 4156 7984 4208
rect 14372 4156 14424 4208
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 6828 4088 6880 4140
rect 4896 4020 4948 4072
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8576 4088 8628 4140
rect 15936 4088 15988 4140
rect 19156 4088 19208 4140
rect 8116 4020 8168 4072
rect 12532 4063 12584 4072
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 13452 4020 13504 4072
rect 7759 3782 7811 3834
rect 7823 3782 7875 3834
rect 7887 3782 7939 3834
rect 7951 3782 8003 3834
rect 14536 3782 14588 3834
rect 14600 3782 14652 3834
rect 14664 3782 14716 3834
rect 14728 3782 14780 3834
rect 7288 3680 7340 3732
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 4370 3238 4422 3290
rect 4434 3238 4486 3290
rect 4498 3238 4550 3290
rect 4562 3238 4614 3290
rect 11148 3238 11200 3290
rect 11212 3238 11264 3290
rect 11276 3238 11328 3290
rect 11340 3238 11392 3290
rect 17925 3238 17977 3290
rect 17989 3238 18041 3290
rect 18053 3238 18105 3290
rect 18117 3238 18169 3290
rect 4252 3000 4304 3052
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 4160 2932 4212 2984
rect 16120 2932 16172 2984
rect 15108 2864 15160 2916
rect 572 2796 624 2848
rect 5080 2796 5132 2848
rect 8300 2796 8352 2848
rect 8668 2796 8720 2848
rect 7759 2694 7811 2746
rect 7823 2694 7875 2746
rect 7887 2694 7939 2746
rect 7951 2694 8003 2746
rect 14536 2694 14588 2746
rect 14600 2694 14652 2746
rect 14664 2694 14716 2746
rect 14728 2694 14780 2746
rect 7656 2524 7708 2576
rect 8300 2456 8352 2508
rect 8944 2524 8996 2576
rect 16948 2524 17000 2576
rect 12256 2456 12308 2508
rect 4370 2150 4422 2202
rect 4434 2150 4486 2202
rect 4498 2150 4550 2202
rect 4562 2150 4614 2202
rect 11148 2150 11200 2202
rect 11212 2150 11264 2202
rect 11276 2150 11328 2202
rect 11340 2150 11392 2202
rect 17925 2150 17977 2202
rect 17989 2150 18041 2202
rect 18053 2150 18105 2202
rect 18117 2150 18169 2202
<< metal2 >>
rect 3330 23933 3386 24733
rect 9586 23933 9642 24733
rect 15842 23933 15898 24733
rect 21914 23933 21970 24733
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 10062 1440 17682
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1780 9994 1808 11086
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1688 8498 1716 8910
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7002 1624 7142
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1780 6798 1808 9930
rect 1872 8974 1900 17614
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 15978 2728 17546
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2424 8906 2452 15914
rect 2792 12102 2820 19071
rect 2976 16658 3004 19926
rect 3344 19378 3372 23933
rect 7733 22332 8029 22352
rect 7789 22330 7813 22332
rect 7869 22330 7893 22332
rect 7949 22330 7973 22332
rect 7811 22278 7813 22330
rect 7875 22278 7887 22330
rect 7949 22278 7951 22330
rect 7789 22276 7813 22278
rect 7869 22276 7893 22278
rect 7949 22276 7973 22278
rect 7733 22256 8029 22276
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 4344 21788 4640 21808
rect 4400 21786 4424 21788
rect 4480 21786 4504 21788
rect 4560 21786 4584 21788
rect 4422 21734 4424 21786
rect 4486 21734 4498 21786
rect 4560 21734 4562 21786
rect 4400 21732 4424 21734
rect 4480 21732 4504 21734
rect 4560 21732 4584 21734
rect 4344 21712 4640 21732
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 4344 20700 4640 20720
rect 4400 20698 4424 20700
rect 4480 20698 4504 20700
rect 4560 20698 4584 20700
rect 4422 20646 4424 20698
rect 4486 20646 4498 20698
rect 4560 20646 4562 20698
rect 4400 20644 4424 20646
rect 4480 20644 4504 20646
rect 4560 20644 4584 20646
rect 4344 20624 4640 20644
rect 4344 19612 4640 19632
rect 4400 19610 4424 19612
rect 4480 19610 4504 19612
rect 4560 19610 4584 19612
rect 4422 19558 4424 19610
rect 4486 19558 4498 19610
rect 4560 19558 4562 19610
rect 4400 19556 4424 19558
rect 4480 19556 4504 19558
rect 4560 19556 4584 19558
rect 4344 19536 4640 19556
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 4344 18524 4640 18544
rect 4400 18522 4424 18524
rect 4480 18522 4504 18524
rect 4560 18522 4584 18524
rect 4422 18470 4424 18522
rect 4486 18470 4498 18522
rect 4560 18470 4562 18522
rect 4400 18468 4424 18470
rect 4480 18468 4504 18470
rect 4560 18468 4584 18470
rect 4344 18448 4640 18468
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15638 2912 15982
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 7954 2452 8842
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2056 6458 2084 6802
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2608 6390 2636 10746
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 10198 2728 10406
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2700 5778 2728 8366
rect 2792 6254 2820 12038
rect 2976 6254 3004 16594
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3528 14618 3556 14894
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 3068 9110 3096 13194
rect 3252 12850 3280 14554
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3436 12866 3464 12922
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3344 12838 3464 12866
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3068 7342 3096 9046
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 3160 4146 3188 11562
rect 3344 5846 3372 12838
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 8430 3556 9522
rect 3620 8634 3648 18090
rect 4344 17436 4640 17456
rect 4400 17434 4424 17436
rect 4480 17434 4504 17436
rect 4560 17434 4584 17436
rect 4422 17382 4424 17434
rect 4486 17382 4498 17434
rect 4560 17382 4562 17434
rect 4400 17380 4424 17382
rect 4480 17380 4504 17382
rect 4560 17380 4584 17382
rect 4344 17360 4640 17380
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7342 3464 7686
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3804 4078 3832 17002
rect 4344 16348 4640 16368
rect 4400 16346 4424 16348
rect 4480 16346 4504 16348
rect 4560 16346 4584 16348
rect 4422 16294 4424 16346
rect 4486 16294 4498 16346
rect 4560 16294 4562 16346
rect 4400 16292 4424 16294
rect 4480 16292 4504 16294
rect 4560 16292 4584 16294
rect 4344 16272 4640 16292
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4344 15260 4640 15280
rect 4400 15258 4424 15260
rect 4480 15258 4504 15260
rect 4560 15258 4584 15260
rect 4422 15206 4424 15258
rect 4486 15206 4498 15258
rect 4560 15206 4562 15258
rect 4400 15204 4424 15206
rect 4480 15204 4504 15206
rect 4560 15204 4584 15206
rect 4344 15184 4640 15204
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 4146 3924 13262
rect 4080 10130 4108 14214
rect 4264 11762 4292 14894
rect 4344 14172 4640 14192
rect 4400 14170 4424 14172
rect 4480 14170 4504 14172
rect 4560 14170 4584 14172
rect 4422 14118 4424 14170
rect 4486 14118 4498 14170
rect 4560 14118 4562 14170
rect 4400 14116 4424 14118
rect 4480 14116 4504 14118
rect 4560 14116 4584 14118
rect 4344 14096 4640 14116
rect 4344 13084 4640 13104
rect 4400 13082 4424 13084
rect 4480 13082 4504 13084
rect 4560 13082 4584 13084
rect 4422 13030 4424 13082
rect 4486 13030 4498 13082
rect 4560 13030 4562 13082
rect 4400 13028 4424 13030
rect 4480 13028 4504 13030
rect 4560 13028 4584 13030
rect 4344 13008 4640 13028
rect 4344 11996 4640 12016
rect 4400 11994 4424 11996
rect 4480 11994 4504 11996
rect 4560 11994 4584 11996
rect 4422 11942 4424 11994
rect 4486 11942 4498 11994
rect 4560 11942 4562 11994
rect 4400 11940 4424 11942
rect 4480 11940 4504 11942
rect 4560 11940 4584 11942
rect 4344 11920 4640 11940
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4344 10908 4640 10928
rect 4400 10906 4424 10908
rect 4480 10906 4504 10908
rect 4560 10906 4584 10908
rect 4422 10854 4424 10906
rect 4486 10854 4498 10906
rect 4560 10854 4562 10906
rect 4400 10852 4424 10854
rect 4480 10852 4504 10854
rect 4560 10852 4584 10854
rect 4344 10832 4640 10852
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4066 9888 4122 9897
rect 4066 9823 4122 9832
rect 4080 9722 4108 9823
rect 4344 9820 4640 9840
rect 4400 9818 4424 9820
rect 4480 9818 4504 9820
rect 4560 9818 4584 9820
rect 4422 9766 4424 9818
rect 4486 9766 4498 9818
rect 4560 9766 4562 9818
rect 4400 9764 4424 9766
rect 4480 9764 4504 9766
rect 4560 9764 4584 9766
rect 4344 9744 4640 9764
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 6866 4016 8910
rect 4068 7948 4120 7954
rect 4172 7936 4200 9590
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4120 7908 4200 7936
rect 4068 7890 4120 7896
rect 4264 7274 4292 8910
rect 4344 8732 4640 8752
rect 4400 8730 4424 8732
rect 4480 8730 4504 8732
rect 4560 8730 4584 8732
rect 4422 8678 4424 8730
rect 4486 8678 4498 8730
rect 4560 8678 4562 8730
rect 4400 8676 4424 8678
rect 4480 8676 4504 8678
rect 4560 8676 4584 8678
rect 4344 8656 4640 8676
rect 4724 8022 4752 10950
rect 4908 10282 4936 15302
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 11354 5028 11766
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4908 10254 5028 10282
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4802 9752 4858 9761
rect 4802 9687 4858 9696
rect 4816 9654 4844 9687
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4344 7644 4640 7664
rect 4400 7642 4424 7644
rect 4480 7642 4504 7644
rect 4560 7642 4584 7644
rect 4422 7590 4424 7642
rect 4486 7590 4498 7642
rect 4560 7590 4562 7642
rect 4400 7588 4424 7590
rect 4480 7588 4504 7590
rect 4560 7588 4584 7590
rect 4344 7568 4640 7588
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4172 5778 4200 6122
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 4172 2990 4200 5714
rect 4264 3058 4292 7210
rect 4344 6556 4640 6576
rect 4400 6554 4424 6556
rect 4480 6554 4504 6556
rect 4560 6554 4584 6556
rect 4422 6502 4424 6554
rect 4486 6502 4498 6554
rect 4560 6502 4562 6554
rect 4400 6500 4424 6502
rect 4480 6500 4504 6502
rect 4560 6500 4584 6502
rect 4344 6480 4640 6500
rect 4344 5468 4640 5488
rect 4400 5466 4424 5468
rect 4480 5466 4504 5468
rect 4560 5466 4584 5468
rect 4422 5414 4424 5466
rect 4486 5414 4498 5466
rect 4560 5414 4562 5466
rect 4400 5412 4424 5414
rect 4480 5412 4504 5414
rect 4560 5412 4584 5414
rect 4344 5392 4640 5412
rect 4908 4826 4936 10066
rect 5000 9450 5028 10254
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5000 7342 5028 9386
rect 5092 9178 5120 15506
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5092 7750 5120 9114
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4344 4380 4640 4400
rect 4400 4378 4424 4380
rect 4480 4378 4504 4380
rect 4560 4378 4584 4380
rect 4422 4326 4424 4378
rect 4486 4326 4498 4378
rect 4560 4326 4562 4378
rect 4400 4324 4424 4326
rect 4480 4324 4504 4326
rect 4560 4324 4584 4326
rect 4344 4304 4640 4324
rect 4908 4078 4936 4762
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4344 3292 4640 3312
rect 4400 3290 4424 3292
rect 4480 3290 4504 3292
rect 4560 3290 4584 3292
rect 4422 3238 4424 3290
rect 4486 3238 4498 3290
rect 4560 3238 4562 3290
rect 4400 3236 4424 3238
rect 4480 3236 4504 3238
rect 4560 3236 4584 3238
rect 4344 3216 4640 3236
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 5092 2854 5120 7686
rect 5184 3058 5212 14350
rect 5276 6322 5304 17070
rect 5368 9761 5396 17138
rect 5354 9752 5410 9761
rect 5354 9687 5410 9696
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5552 7206 5580 9046
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 6380 4826 6408 20946
rect 7392 19174 7420 21898
rect 7733 21244 8029 21264
rect 7789 21242 7813 21244
rect 7869 21242 7893 21244
rect 7949 21242 7973 21244
rect 7811 21190 7813 21242
rect 7875 21190 7887 21242
rect 7949 21190 7951 21242
rect 7789 21188 7813 21190
rect 7869 21188 7893 21190
rect 7949 21188 7973 21190
rect 7733 21168 8029 21188
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 7733 20156 8029 20176
rect 7789 20154 7813 20156
rect 7869 20154 7893 20156
rect 7949 20154 7973 20156
rect 7811 20102 7813 20154
rect 7875 20102 7887 20154
rect 7949 20102 7951 20154
rect 7789 20100 7813 20102
rect 7869 20100 7893 20102
rect 7949 20100 7973 20102
rect 7733 20080 8029 20100
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6748 16250 6776 17070
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6748 15910 6776 16186
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6932 13394 6960 18022
rect 7392 16046 7420 19110
rect 7733 19068 8029 19088
rect 7789 19066 7813 19068
rect 7869 19066 7893 19068
rect 7949 19066 7973 19068
rect 7811 19014 7813 19066
rect 7875 19014 7887 19066
rect 7949 19014 7951 19066
rect 7789 19012 7813 19014
rect 7869 19012 7893 19014
rect 7949 19012 7973 19014
rect 7733 18992 8029 19012
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6932 12986 6960 13330
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6748 9926 6776 11222
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6840 9654 6868 11222
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6564 7342 6592 9590
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7024 9042 7052 9318
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8430 7052 8978
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 7002 6592 7278
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6564 4690 6592 6938
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 584 800 612 2790
rect 4344 2204 4640 2224
rect 4400 2202 4424 2204
rect 4480 2202 4504 2204
rect 4560 2202 4584 2204
rect 4422 2150 4424 2202
rect 4486 2150 4498 2202
rect 4560 2150 4562 2202
rect 4400 2148 4424 2150
rect 4480 2148 4504 2150
rect 4560 2148 4584 2150
rect 4344 2128 4640 2148
rect 6656 800 6684 7142
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6840 6390 6868 6870
rect 7024 6798 7052 8366
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6840 4146 6868 6326
rect 7116 4690 7144 15982
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7300 3738 7328 8366
rect 7576 4690 7604 18090
rect 7733 17980 8029 18000
rect 7789 17978 7813 17980
rect 7869 17978 7893 17980
rect 7949 17978 7973 17980
rect 7811 17926 7813 17978
rect 7875 17926 7887 17978
rect 7949 17926 7951 17978
rect 7789 17924 7813 17926
rect 7869 17924 7893 17926
rect 7949 17924 7973 17926
rect 7733 17904 8029 17924
rect 7733 16892 8029 16912
rect 7789 16890 7813 16892
rect 7869 16890 7893 16892
rect 7949 16890 7973 16892
rect 7811 16838 7813 16890
rect 7875 16838 7887 16890
rect 7949 16838 7951 16890
rect 7789 16836 7813 16838
rect 7869 16836 7893 16838
rect 7949 16836 7973 16838
rect 7733 16816 8029 16836
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 11354 7696 15982
rect 7733 15804 8029 15824
rect 7789 15802 7813 15804
rect 7869 15802 7893 15804
rect 7949 15802 7973 15804
rect 7811 15750 7813 15802
rect 7875 15750 7887 15802
rect 7949 15750 7951 15802
rect 7789 15748 7813 15750
rect 7869 15748 7893 15750
rect 7949 15748 7973 15750
rect 7733 15728 8029 15748
rect 7733 14716 8029 14736
rect 7789 14714 7813 14716
rect 7869 14714 7893 14716
rect 7949 14714 7973 14716
rect 7811 14662 7813 14714
rect 7875 14662 7887 14714
rect 7949 14662 7951 14714
rect 7789 14660 7813 14662
rect 7869 14660 7893 14662
rect 7949 14660 7973 14662
rect 7733 14640 8029 14660
rect 7733 13628 8029 13648
rect 7789 13626 7813 13628
rect 7869 13626 7893 13628
rect 7949 13626 7973 13628
rect 7811 13574 7813 13626
rect 7875 13574 7887 13626
rect 7949 13574 7951 13626
rect 7789 13572 7813 13574
rect 7869 13572 7893 13574
rect 7949 13572 7973 13574
rect 7733 13552 8029 13572
rect 7733 12540 8029 12560
rect 7789 12538 7813 12540
rect 7869 12538 7893 12540
rect 7949 12538 7973 12540
rect 7811 12486 7813 12538
rect 7875 12486 7887 12538
rect 7949 12486 7951 12538
rect 7789 12484 7813 12486
rect 7869 12484 7893 12486
rect 7949 12484 7973 12486
rect 7733 12464 8029 12484
rect 7733 11452 8029 11472
rect 7789 11450 7813 11452
rect 7869 11450 7893 11452
rect 7949 11450 7973 11452
rect 7811 11398 7813 11450
rect 7875 11398 7887 11450
rect 7949 11398 7951 11450
rect 7789 11396 7813 11398
rect 7869 11396 7893 11398
rect 7949 11396 7973 11398
rect 7733 11376 8029 11396
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7733 10364 8029 10384
rect 7789 10362 7813 10364
rect 7869 10362 7893 10364
rect 7949 10362 7973 10364
rect 7811 10310 7813 10362
rect 7875 10310 7887 10362
rect 7949 10310 7951 10362
rect 7789 10308 7813 10310
rect 7869 10308 7893 10310
rect 7949 10308 7973 10310
rect 7733 10288 8029 10308
rect 7733 9276 8029 9296
rect 7789 9274 7813 9276
rect 7869 9274 7893 9276
rect 7949 9274 7973 9276
rect 7811 9222 7813 9274
rect 7875 9222 7887 9274
rect 7949 9222 7951 9274
rect 7789 9220 7813 9222
rect 7869 9220 7893 9222
rect 7949 9220 7973 9222
rect 7733 9200 8029 9220
rect 7733 8188 8029 8208
rect 7789 8186 7813 8188
rect 7869 8186 7893 8188
rect 7949 8186 7973 8188
rect 7811 8134 7813 8186
rect 7875 8134 7887 8186
rect 7949 8134 7951 8186
rect 7789 8132 7813 8134
rect 7869 8132 7893 8134
rect 7949 8132 7973 8134
rect 7733 8112 8029 8132
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7668 4282 7696 7754
rect 7733 7100 8029 7120
rect 7789 7098 7813 7100
rect 7869 7098 7893 7100
rect 7949 7098 7973 7100
rect 7811 7046 7813 7098
rect 7875 7046 7887 7098
rect 7949 7046 7951 7098
rect 7789 7044 7813 7046
rect 7869 7044 7893 7046
rect 7949 7044 7973 7046
rect 7733 7024 8029 7044
rect 7733 6012 8029 6032
rect 7789 6010 7813 6012
rect 7869 6010 7893 6012
rect 7949 6010 7973 6012
rect 7811 5958 7813 6010
rect 7875 5958 7887 6010
rect 7949 5958 7951 6010
rect 7789 5956 7813 5958
rect 7869 5956 7893 5958
rect 7949 5956 7973 5958
rect 7733 5936 8029 5956
rect 7733 4924 8029 4944
rect 7789 4922 7813 4924
rect 7869 4922 7893 4924
rect 7949 4922 7973 4924
rect 7811 4870 7813 4922
rect 7875 4870 7887 4922
rect 7949 4870 7951 4922
rect 7789 4868 7813 4870
rect 7869 4868 7893 4870
rect 7949 4868 7973 4870
rect 7733 4848 8029 4868
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7668 2582 7696 4218
rect 7944 4214 7972 4558
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 4078 7972 4150
rect 8128 4078 8156 19246
rect 8312 15978 8340 20810
rect 8392 20324 8444 20330
rect 8392 20266 8444 20272
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8404 8566 8432 20266
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8496 14618 8524 19110
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10674 8524 10950
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8404 4758 8432 8502
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8588 4146 8616 22102
rect 9220 21412 9272 21418
rect 9220 21354 9272 21360
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 11694 8708 19314
rect 8864 19174 8892 19926
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8772 11370 8800 12174
rect 8680 11342 8800 11370
rect 8680 10538 8708 11342
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8772 10538 8800 11222
rect 8864 11014 8892 19110
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9048 12306 9076 14554
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9140 11898 9168 12582
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7733 3836 8029 3856
rect 7789 3834 7813 3836
rect 7869 3834 7893 3836
rect 7949 3834 7973 3836
rect 7811 3782 7813 3834
rect 7875 3782 7887 3834
rect 7949 3782 7951 3834
rect 7789 3780 7813 3782
rect 7869 3780 7893 3782
rect 7949 3780 7973 3782
rect 7733 3760 8029 3780
rect 8680 2854 8708 10474
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 7733 2748 8029 2768
rect 7789 2746 7813 2748
rect 7869 2746 7893 2748
rect 7949 2746 7973 2748
rect 7811 2694 7813 2746
rect 7875 2694 7887 2746
rect 7949 2694 7951 2746
rect 7789 2692 7813 2694
rect 7869 2692 7893 2694
rect 7949 2692 7973 2694
rect 7733 2672 8029 2692
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8312 2514 8340 2790
rect 8956 2582 8984 11086
rect 9048 9518 9076 11494
rect 9128 10464 9180 10470
rect 9232 10418 9260 21354
rect 9600 20602 9628 23933
rect 14510 22332 14806 22352
rect 14566 22330 14590 22332
rect 14646 22330 14670 22332
rect 14726 22330 14750 22332
rect 14588 22278 14590 22330
rect 14652 22278 14664 22330
rect 14726 22278 14728 22330
rect 14566 22276 14590 22278
rect 14646 22276 14670 22278
rect 14726 22276 14750 22278
rect 14510 22256 14806 22276
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 11122 21788 11418 21808
rect 11178 21786 11202 21788
rect 11258 21786 11282 21788
rect 11338 21786 11362 21788
rect 11200 21734 11202 21786
rect 11264 21734 11276 21786
rect 11338 21734 11340 21786
rect 11178 21732 11202 21734
rect 11258 21732 11282 21734
rect 11338 21732 11362 21734
rect 11122 21712 11418 21732
rect 12072 21616 12124 21622
rect 12072 21558 12124 21564
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 11762 9536 16934
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11506 9536 11698
rect 9600 11558 9628 14418
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 11694 9720 14214
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9416 11478 9536 11506
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9416 11286 9444 11478
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10418 9352 10474
rect 9180 10412 9352 10418
rect 9128 10406 9352 10412
rect 9140 10390 9352 10406
rect 9508 9654 9536 11290
rect 9692 10470 9720 11630
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9232 6798 9260 9590
rect 9600 9042 9628 9658
rect 9876 9654 9904 11086
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9876 9382 9904 9590
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9968 9042 9996 15846
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10060 10010 10088 14554
rect 10152 10198 10180 19994
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11558 10364 11630
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10060 9982 10180 10010
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 9722 10088 9862
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9600 8634 9628 8978
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 6916 9444 7754
rect 9588 6928 9640 6934
rect 9416 6888 9588 6916
rect 9588 6870 9640 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 10152 5642 10180 9982
rect 10428 6866 10456 17682
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10704 3602 10732 20878
rect 11122 20700 11418 20720
rect 11178 20698 11202 20700
rect 11258 20698 11282 20700
rect 11338 20698 11362 20700
rect 11200 20646 11202 20698
rect 11264 20646 11276 20698
rect 11338 20646 11340 20698
rect 11178 20644 11202 20646
rect 11258 20644 11282 20646
rect 11338 20644 11362 20646
rect 11122 20624 11418 20644
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11122 19612 11418 19632
rect 11178 19610 11202 19612
rect 11258 19610 11282 19612
rect 11338 19610 11362 19612
rect 11200 19558 11202 19610
rect 11264 19558 11276 19610
rect 11338 19558 11340 19610
rect 11178 19556 11202 19558
rect 11258 19556 11282 19558
rect 11338 19556 11362 19558
rect 11122 19536 11418 19556
rect 11122 18524 11418 18544
rect 11178 18522 11202 18524
rect 11258 18522 11282 18524
rect 11338 18522 11362 18524
rect 11200 18470 11202 18522
rect 11264 18470 11276 18522
rect 11338 18470 11340 18522
rect 11178 18468 11202 18470
rect 11258 18468 11282 18470
rect 11338 18468 11362 18470
rect 11122 18448 11418 18468
rect 11122 17436 11418 17456
rect 11178 17434 11202 17436
rect 11258 17434 11282 17436
rect 11338 17434 11362 17436
rect 11200 17382 11202 17434
rect 11264 17382 11276 17434
rect 11338 17382 11340 17434
rect 11178 17380 11202 17382
rect 11258 17380 11282 17382
rect 11338 17380 11362 17382
rect 11122 17360 11418 17380
rect 11122 16348 11418 16368
rect 11178 16346 11202 16348
rect 11258 16346 11282 16348
rect 11338 16346 11362 16348
rect 11200 16294 11202 16346
rect 11264 16294 11276 16346
rect 11338 16294 11340 16346
rect 11178 16292 11202 16294
rect 11258 16292 11282 16294
rect 11338 16292 11362 16294
rect 11122 16272 11418 16292
rect 11122 15260 11418 15280
rect 11178 15258 11202 15260
rect 11258 15258 11282 15260
rect 11338 15258 11362 15260
rect 11200 15206 11202 15258
rect 11264 15206 11276 15258
rect 11338 15206 11340 15258
rect 11178 15204 11202 15206
rect 11258 15204 11282 15206
rect 11338 15204 11362 15206
rect 11122 15184 11418 15204
rect 11532 15026 11560 19858
rect 11796 19848 11848 19854
rect 11992 19802 12020 21490
rect 11848 19796 12020 19802
rect 11796 19790 12020 19796
rect 11808 19774 12020 19790
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11122 14172 11418 14192
rect 11178 14170 11202 14172
rect 11258 14170 11282 14172
rect 11338 14170 11362 14172
rect 11200 14118 11202 14170
rect 11264 14118 11276 14170
rect 11338 14118 11340 14170
rect 11178 14116 11202 14118
rect 11258 14116 11282 14118
rect 11338 14116 11362 14118
rect 11122 14096 11418 14116
rect 11122 13084 11418 13104
rect 11178 13082 11202 13084
rect 11258 13082 11282 13084
rect 11338 13082 11362 13084
rect 11200 13030 11202 13082
rect 11264 13030 11276 13082
rect 11338 13030 11340 13082
rect 11178 13028 11202 13030
rect 11258 13028 11282 13030
rect 11338 13028 11362 13030
rect 11122 13008 11418 13028
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11354 10916 12038
rect 11122 11996 11418 12016
rect 11178 11994 11202 11996
rect 11258 11994 11282 11996
rect 11338 11994 11362 11996
rect 11200 11942 11202 11994
rect 11264 11942 11276 11994
rect 11338 11942 11340 11994
rect 11178 11940 11202 11942
rect 11258 11940 11282 11942
rect 11338 11940 11362 11942
rect 11122 11920 11418 11940
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11122 10908 11418 10928
rect 11178 10906 11202 10908
rect 11258 10906 11282 10908
rect 11338 10906 11362 10908
rect 11200 10854 11202 10906
rect 11264 10854 11276 10906
rect 11338 10854 11340 10906
rect 11178 10852 11202 10854
rect 11258 10852 11282 10854
rect 11338 10852 11362 10854
rect 11122 10832 11418 10852
rect 11532 10742 11560 10950
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11122 9820 11418 9840
rect 11178 9818 11202 9820
rect 11258 9818 11282 9820
rect 11338 9818 11362 9820
rect 11200 9766 11202 9818
rect 11264 9766 11276 9818
rect 11338 9766 11340 9818
rect 11178 9764 11202 9766
rect 11258 9764 11282 9766
rect 11338 9764 11362 9766
rect 11122 9744 11418 9764
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11122 8732 11418 8752
rect 11178 8730 11202 8732
rect 11258 8730 11282 8732
rect 11338 8730 11362 8732
rect 11200 8678 11202 8730
rect 11264 8678 11276 8730
rect 11338 8678 11340 8730
rect 11178 8676 11202 8678
rect 11258 8676 11282 8678
rect 11338 8676 11362 8678
rect 11122 8656 11418 8676
rect 11532 8566 11560 8978
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11122 7644 11418 7664
rect 11178 7642 11202 7644
rect 11258 7642 11282 7644
rect 11338 7642 11362 7644
rect 11200 7590 11202 7642
rect 11264 7590 11276 7642
rect 11338 7590 11340 7642
rect 11178 7588 11202 7590
rect 11258 7588 11282 7590
rect 11338 7588 11362 7590
rect 11122 7568 11418 7588
rect 11532 7546 11560 8502
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11122 6556 11418 6576
rect 11178 6554 11202 6556
rect 11258 6554 11282 6556
rect 11338 6554 11362 6556
rect 11200 6502 11202 6554
rect 11264 6502 11276 6554
rect 11338 6502 11340 6554
rect 11178 6500 11202 6502
rect 11258 6500 11282 6502
rect 11338 6500 11362 6502
rect 11122 6480 11418 6500
rect 11532 5710 11560 6598
rect 11624 5914 11652 17614
rect 11716 16726 11744 18226
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 12646 11744 16662
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11716 11218 11744 12106
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11716 6662 11744 7958
rect 11808 7410 11836 12718
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11900 9518 11928 11834
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11992 8022 12020 19774
rect 12084 12102 12112 21558
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12728 20602 12756 20946
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12176 17814 12204 20538
rect 12728 20466 12756 20538
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11082 12112 12038
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 12084 5642 12112 11018
rect 12176 5778 12204 17750
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13096 16658 13124 17138
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 12322 12480 14758
rect 12452 12294 12664 12322
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12268 11762 12296 11834
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12544 11626 12572 12174
rect 12348 11620 12400 11626
rect 12532 11620 12584 11626
rect 12400 11580 12480 11608
rect 12348 11562 12400 11568
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11122 5468 11418 5488
rect 11178 5466 11202 5468
rect 11258 5466 11282 5468
rect 11338 5466 11362 5468
rect 11200 5414 11202 5466
rect 11264 5414 11276 5466
rect 11338 5414 11340 5466
rect 11178 5412 11202 5414
rect 11258 5412 11282 5414
rect 11338 5412 11362 5414
rect 11122 5392 11418 5412
rect 11122 4380 11418 4400
rect 11178 4378 11202 4380
rect 11258 4378 11282 4380
rect 11338 4378 11362 4380
rect 11200 4326 11202 4378
rect 11264 4326 11276 4378
rect 11338 4326 11340 4378
rect 11178 4324 11202 4326
rect 11258 4324 11282 4326
rect 11338 4324 11362 4326
rect 11122 4304 11418 4324
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 11122 3292 11418 3312
rect 11178 3290 11202 3292
rect 11258 3290 11282 3292
rect 11338 3290 11362 3292
rect 11200 3238 11202 3290
rect 11264 3238 11276 3290
rect 11338 3238 11340 3290
rect 11178 3236 11202 3238
rect 11258 3236 11282 3238
rect 11338 3236 11362 3238
rect 11122 3216 11418 3236
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 12268 2514 12296 10406
rect 12452 7546 12480 11580
rect 12532 11562 12584 11568
rect 12636 9659 12664 12294
rect 13004 11898 13032 16594
rect 13096 14550 13124 16594
rect 13188 15026 13216 21422
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18834 13400 19246
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12728 11694 12756 11834
rect 13188 11762 13216 14962
rect 13280 14414 13308 18158
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12622 9650 12678 9659
rect 12622 9585 12678 9594
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 9382 12572 9454
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12360 6730 12388 7210
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12544 4078 12572 9318
rect 12728 4078 12756 10542
rect 12820 7954 12848 11562
rect 13188 11286 13216 11562
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 9654 12940 10542
rect 13280 9761 13308 14350
rect 13464 13274 13492 21830
rect 14510 21244 14806 21264
rect 14566 21242 14590 21244
rect 14646 21242 14670 21244
rect 14726 21242 14750 21244
rect 14588 21190 14590 21242
rect 14652 21190 14664 21242
rect 14726 21190 14728 21242
rect 14566 21188 14590 21190
rect 14646 21188 14670 21190
rect 14726 21188 14750 21190
rect 14510 21168 14806 21188
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14510 20156 14806 20176
rect 14566 20154 14590 20156
rect 14646 20154 14670 20156
rect 14726 20154 14750 20156
rect 14588 20102 14590 20154
rect 14652 20102 14664 20154
rect 14726 20102 14728 20154
rect 14566 20100 14590 20102
rect 14646 20100 14670 20102
rect 14726 20100 14750 20102
rect 14510 20080 14806 20100
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13648 15858 13676 19246
rect 14510 19068 14806 19088
rect 14566 19066 14590 19068
rect 14646 19066 14670 19068
rect 14726 19066 14750 19068
rect 14588 19014 14590 19066
rect 14652 19014 14664 19066
rect 14726 19014 14728 19066
rect 14566 19012 14590 19014
rect 14646 19012 14670 19014
rect 14726 19012 14750 19014
rect 14510 18992 14806 19012
rect 14510 17980 14806 18000
rect 14566 17978 14590 17980
rect 14646 17978 14670 17980
rect 14726 17978 14750 17980
rect 14588 17926 14590 17978
rect 14652 17926 14664 17978
rect 14726 17926 14728 17978
rect 14566 17924 14590 17926
rect 14646 17924 14670 17926
rect 14726 17924 14750 17926
rect 14510 17904 14806 17924
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13372 13246 13492 13274
rect 13556 15830 13676 15858
rect 13372 12730 13400 13246
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 12918 13492 13126
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13372 12702 13492 12730
rect 13266 9752 13322 9761
rect 13266 9687 13322 9696
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 12898 8528 12954 8537
rect 12898 8463 12900 8472
rect 12952 8463 12954 8472
rect 12900 8434 12952 8440
rect 13004 8378 13032 9551
rect 12912 8350 13032 8378
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12912 7342 12940 8350
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 11122 2204 11418 2224
rect 11178 2202 11202 2204
rect 11258 2202 11282 2204
rect 11338 2202 11362 2204
rect 11200 2150 11202 2202
rect 11264 2150 11276 2202
rect 11338 2150 11340 2202
rect 11178 2148 11202 2150
rect 11258 2148 11282 2150
rect 11338 2148 11362 2150
rect 11122 2128 11418 2148
rect 12912 800 12940 7278
rect 13464 4078 13492 12702
rect 13556 9178 13584 15830
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12986 13676 13262
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 12866 13768 15574
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13648 12838 13768 12866
rect 13648 11626 13676 12838
rect 13832 12306 13860 14758
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13924 10674 13952 14894
rect 14016 12730 14044 16730
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 12918 14136 14826
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14016 12702 14136 12730
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13740 4622 13768 9590
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9110 13860 9454
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13924 7478 13952 9590
rect 14016 9194 14044 12582
rect 14108 10130 14136 12702
rect 14200 10266 14228 15982
rect 14292 15026 14320 16186
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14384 12866 14412 17750
rect 14510 16892 14806 16912
rect 14566 16890 14590 16892
rect 14646 16890 14670 16892
rect 14726 16890 14750 16892
rect 14588 16838 14590 16890
rect 14652 16838 14664 16890
rect 14726 16838 14728 16890
rect 14566 16836 14590 16838
rect 14646 16836 14670 16838
rect 14726 16836 14750 16838
rect 14510 16816 14806 16836
rect 14510 15804 14806 15824
rect 14566 15802 14590 15804
rect 14646 15802 14670 15804
rect 14726 15802 14750 15804
rect 14588 15750 14590 15802
rect 14652 15750 14664 15802
rect 14726 15750 14728 15802
rect 14566 15748 14590 15750
rect 14646 15748 14670 15750
rect 14726 15748 14750 15750
rect 14510 15728 14806 15748
rect 14510 14716 14806 14736
rect 14566 14714 14590 14716
rect 14646 14714 14670 14716
rect 14726 14714 14750 14716
rect 14588 14662 14590 14714
rect 14652 14662 14664 14714
rect 14726 14662 14728 14714
rect 14566 14660 14590 14662
rect 14646 14660 14670 14662
rect 14726 14660 14750 14662
rect 14510 14640 14806 14660
rect 14510 13628 14806 13648
rect 14566 13626 14590 13628
rect 14646 13626 14670 13628
rect 14726 13626 14750 13628
rect 14588 13574 14590 13626
rect 14652 13574 14664 13626
rect 14726 13574 14728 13626
rect 14566 13572 14590 13574
rect 14646 13572 14670 13574
rect 14726 13572 14750 13574
rect 14510 13552 14806 13572
rect 14292 12838 14412 12866
rect 14292 12782 14320 12838
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14292 9518 14320 12582
rect 14384 10742 14412 12650
rect 14510 12540 14806 12560
rect 14566 12538 14590 12540
rect 14646 12538 14670 12540
rect 14726 12538 14750 12540
rect 14588 12486 14590 12538
rect 14652 12486 14664 12538
rect 14726 12486 14728 12538
rect 14566 12484 14590 12486
rect 14646 12484 14670 12486
rect 14726 12484 14750 12486
rect 14510 12464 14806 12484
rect 14510 11452 14806 11472
rect 14566 11450 14590 11452
rect 14646 11450 14670 11452
rect 14726 11450 14750 11452
rect 14588 11398 14590 11450
rect 14652 11398 14664 11450
rect 14726 11398 14728 11450
rect 14566 11396 14590 11398
rect 14646 11396 14670 11398
rect 14726 11396 14750 11398
rect 14510 11376 14806 11396
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14016 9166 14136 9194
rect 14108 9110 14136 9166
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8362 14136 9046
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 14108 6186 14136 8298
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 14384 4214 14412 10678
rect 14510 10364 14806 10384
rect 14566 10362 14590 10364
rect 14646 10362 14670 10364
rect 14726 10362 14750 10364
rect 14588 10310 14590 10362
rect 14652 10310 14664 10362
rect 14726 10310 14728 10362
rect 14566 10308 14590 10310
rect 14646 10308 14670 10310
rect 14726 10308 14750 10310
rect 14510 10288 14806 10308
rect 14510 9276 14806 9296
rect 14566 9274 14590 9276
rect 14646 9274 14670 9276
rect 14726 9274 14750 9276
rect 14588 9222 14590 9274
rect 14652 9222 14664 9274
rect 14726 9222 14728 9274
rect 14566 9220 14590 9222
rect 14646 9220 14670 9222
rect 14726 9220 14750 9222
rect 14510 9200 14806 9220
rect 14844 9042 14872 20334
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14936 10130 14964 12854
rect 15028 12714 15056 19654
rect 15120 12782 15148 20198
rect 15304 17066 15332 22034
rect 15856 20330 15884 23933
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 17899 21788 18195 21808
rect 17955 21786 17979 21788
rect 18035 21786 18059 21788
rect 18115 21786 18139 21788
rect 17977 21734 17979 21786
rect 18041 21734 18053 21786
rect 18115 21734 18117 21786
rect 17955 21732 17979 21734
rect 18035 21732 18059 21734
rect 18115 21732 18139 21734
rect 17899 21712 18195 21732
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16304 21412 16356 21418
rect 16304 21354 16356 21360
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 15570 15332 17002
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14510 8188 14806 8208
rect 14566 8186 14590 8188
rect 14646 8186 14670 8188
rect 14726 8186 14750 8188
rect 14588 8134 14590 8186
rect 14652 8134 14664 8186
rect 14726 8134 14728 8186
rect 14566 8132 14590 8134
rect 14646 8132 14670 8134
rect 14726 8132 14750 8134
rect 14510 8112 14806 8132
rect 14510 7100 14806 7120
rect 14566 7098 14590 7100
rect 14646 7098 14670 7100
rect 14726 7098 14750 7100
rect 14588 7046 14590 7098
rect 14652 7046 14664 7098
rect 14726 7046 14728 7098
rect 14566 7044 14590 7046
rect 14646 7044 14670 7046
rect 14726 7044 14750 7046
rect 14510 7024 14806 7044
rect 14936 6934 14964 10066
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15028 8634 15056 8774
rect 15120 8634 15148 12718
rect 15212 11014 15240 15302
rect 15396 13190 15424 17478
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15672 12322 15700 17546
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15580 12294 15700 12322
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14510 6012 14806 6032
rect 14566 6010 14590 6012
rect 14646 6010 14670 6012
rect 14726 6010 14750 6012
rect 14588 5958 14590 6010
rect 14652 5958 14664 6010
rect 14726 5958 14728 6010
rect 14566 5956 14590 5958
rect 14646 5956 14670 5958
rect 14726 5956 14750 5958
rect 14510 5936 14806 5956
rect 14510 4924 14806 4944
rect 14566 4922 14590 4924
rect 14646 4922 14670 4924
rect 14726 4922 14750 4924
rect 14588 4870 14590 4922
rect 14652 4870 14664 4922
rect 14726 4870 14728 4922
rect 14566 4868 14590 4870
rect 14646 4868 14670 4870
rect 14726 4868 14750 4870
rect 14510 4848 14806 4868
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 14510 3836 14806 3856
rect 14566 3834 14590 3836
rect 14646 3834 14670 3836
rect 14726 3834 14750 3836
rect 14588 3782 14590 3834
rect 14652 3782 14664 3834
rect 14726 3782 14728 3834
rect 14566 3780 14590 3782
rect 14646 3780 14670 3782
rect 14726 3780 14750 3782
rect 14510 3760 14806 3780
rect 15120 2922 15148 8570
rect 15212 7274 15240 10950
rect 15580 9654 15608 12294
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15304 8430 15332 9386
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15488 8430 15516 8570
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15672 7410 15700 10474
rect 15856 10266 15884 14826
rect 16316 13274 16344 21354
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16408 19922 16436 20946
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16408 16998 16436 19858
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16500 13394 16528 19178
rect 16592 16726 16620 21286
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16684 19922 16712 20878
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16316 13246 16528 13274
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15842 9616 15898 9625
rect 15842 9551 15898 9560
rect 15750 8528 15806 8537
rect 15750 8463 15752 8472
rect 15804 8463 15806 8472
rect 15752 8434 15804 8440
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6390 15332 6802
rect 15672 6798 15700 7346
rect 15856 6934 15884 9551
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15764 6322 15792 6598
rect 15856 6458 15884 6734
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15948 4146 15976 11562
rect 16132 8838 16160 11630
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16132 2990 16160 8774
rect 16316 6730 16344 9862
rect 16408 6798 16436 10542
rect 16500 9926 16528 13246
rect 16592 11558 16620 16526
rect 16684 12238 16712 19858
rect 16776 16590 16804 21014
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16868 16726 16896 18702
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16960 13462 16988 21422
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 17338 17080 20198
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17052 14482 17080 17274
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16776 12170 16804 13398
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 10062 16620 11494
rect 17144 10606 17172 13330
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16592 9518 16620 9998
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16868 4826 16896 7890
rect 16960 7818 16988 9998
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14510 2748 14806 2768
rect 14566 2746 14590 2748
rect 14646 2746 14670 2748
rect 14726 2746 14750 2748
rect 14588 2694 14590 2746
rect 14652 2694 14664 2746
rect 14726 2694 14728 2746
rect 14566 2692 14590 2694
rect 14646 2692 14670 2694
rect 14726 2692 14750 2694
rect 14510 2672 14806 2692
rect 16960 2582 16988 7754
rect 17236 5370 17264 18838
rect 17328 14414 17356 18906
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17328 6254 17356 13466
rect 17420 10674 17448 20810
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17512 13530 17540 20334
rect 17604 19854 17632 21082
rect 17899 20700 18195 20720
rect 17955 20698 17979 20700
rect 18035 20698 18059 20700
rect 18115 20698 18139 20700
rect 17977 20646 17979 20698
rect 18041 20646 18053 20698
rect 18115 20646 18117 20698
rect 17955 20644 17979 20646
rect 18035 20644 18059 20646
rect 18115 20644 18139 20646
rect 17899 20624 18195 20644
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17604 18902 17632 19790
rect 17899 19612 18195 19632
rect 17955 19610 17979 19612
rect 18035 19610 18059 19612
rect 18115 19610 18139 19612
rect 17977 19558 17979 19610
rect 18041 19558 18053 19610
rect 18115 19558 18117 19610
rect 17955 19556 17979 19558
rect 18035 19556 18059 19558
rect 18115 19556 18139 19558
rect 17899 19536 18195 19556
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17899 18524 18195 18544
rect 17955 18522 17979 18524
rect 18035 18522 18059 18524
rect 18115 18522 18139 18524
rect 17977 18470 17979 18522
rect 18041 18470 18053 18522
rect 18115 18470 18117 18522
rect 17955 18468 17979 18470
rect 18035 18468 18059 18470
rect 18115 18468 18139 18470
rect 17899 18448 18195 18468
rect 18984 18222 19012 21558
rect 19720 21486 19748 21898
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19904 21146 19932 21422
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 17899 17436 18195 17456
rect 17955 17434 17979 17436
rect 18035 17434 18059 17436
rect 18115 17434 18139 17436
rect 17977 17382 17979 17434
rect 18041 17382 18053 17434
rect 18115 17382 18117 17434
rect 17955 17380 17979 17382
rect 18035 17380 18059 17382
rect 18115 17380 18139 17382
rect 17899 17360 18195 17380
rect 17899 16348 18195 16368
rect 17955 16346 17979 16348
rect 18035 16346 18059 16348
rect 18115 16346 18139 16348
rect 17977 16294 17979 16346
rect 18041 16294 18053 16346
rect 18115 16294 18117 16346
rect 17955 16292 17979 16294
rect 18035 16292 18059 16294
rect 18115 16292 18139 16294
rect 17899 16272 18195 16292
rect 17899 15260 18195 15280
rect 17955 15258 17979 15260
rect 18035 15258 18059 15260
rect 18115 15258 18139 15260
rect 17977 15206 17979 15258
rect 18041 15206 18053 15258
rect 18115 15206 18117 15258
rect 17955 15204 17979 15206
rect 18035 15204 18059 15206
rect 18115 15204 18139 15206
rect 17899 15184 18195 15204
rect 19246 14784 19302 14793
rect 19246 14719 19302 14728
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17788 6866 17816 14350
rect 17899 14172 18195 14192
rect 17955 14170 17979 14172
rect 18035 14170 18059 14172
rect 18115 14170 18139 14172
rect 17977 14118 17979 14170
rect 18041 14118 18053 14170
rect 18115 14118 18117 14170
rect 17955 14116 17979 14118
rect 18035 14116 18059 14118
rect 18115 14116 18139 14118
rect 17899 14096 18195 14116
rect 17899 13084 18195 13104
rect 17955 13082 17979 13084
rect 18035 13082 18059 13084
rect 18115 13082 18139 13084
rect 17977 13030 17979 13082
rect 18041 13030 18053 13082
rect 18115 13030 18117 13082
rect 17955 13028 17979 13030
rect 18035 13028 18059 13030
rect 18115 13028 18139 13030
rect 17899 13008 18195 13028
rect 17899 11996 18195 12016
rect 17955 11994 17979 11996
rect 18035 11994 18059 11996
rect 18115 11994 18139 11996
rect 17977 11942 17979 11994
rect 18041 11942 18053 11994
rect 18115 11942 18117 11994
rect 17955 11940 17979 11942
rect 18035 11940 18059 11942
rect 18115 11940 18139 11942
rect 17899 11920 18195 11940
rect 17899 10908 18195 10928
rect 17955 10906 17979 10908
rect 18035 10906 18059 10908
rect 18115 10906 18139 10908
rect 17977 10854 17979 10906
rect 18041 10854 18053 10906
rect 18115 10854 18117 10906
rect 17955 10852 17979 10854
rect 18035 10852 18059 10854
rect 18115 10852 18139 10854
rect 17899 10832 18195 10852
rect 18248 10538 18276 14418
rect 19260 12850 19288 14719
rect 19352 14618 19380 20198
rect 20272 18086 20300 21014
rect 21928 19990 21956 23933
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18340 10470 18368 11766
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 17899 9820 18195 9840
rect 17955 9818 17979 9820
rect 18035 9818 18059 9820
rect 18115 9818 18139 9820
rect 17977 9766 17979 9818
rect 18041 9766 18053 9818
rect 18115 9766 18117 9818
rect 17955 9764 17979 9766
rect 18035 9764 18059 9766
rect 18115 9764 18139 9766
rect 17899 9744 18195 9764
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 17899 8732 18195 8752
rect 17955 8730 17979 8732
rect 18035 8730 18059 8732
rect 18115 8730 18139 8732
rect 17977 8678 17979 8730
rect 18041 8678 18053 8730
rect 18115 8678 18117 8730
rect 17955 8676 17979 8678
rect 18035 8676 18059 8678
rect 18115 8676 18139 8678
rect 17899 8656 18195 8676
rect 17899 7644 18195 7664
rect 17955 7642 17979 7644
rect 18035 7642 18059 7644
rect 18115 7642 18139 7644
rect 17977 7590 17979 7642
rect 18041 7590 18053 7642
rect 18115 7590 18117 7642
rect 17955 7588 17979 7590
rect 18035 7588 18059 7590
rect 18115 7588 18139 7590
rect 17899 7568 18195 7588
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 18248 6662 18276 9658
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 17899 6556 18195 6576
rect 17955 6554 17979 6556
rect 18035 6554 18059 6556
rect 18115 6554 18139 6556
rect 17977 6502 17979 6554
rect 18041 6502 18053 6554
rect 18115 6502 18117 6554
rect 17955 6500 17979 6502
rect 18035 6500 18059 6502
rect 18115 6500 18139 6502
rect 17899 6480 18195 6500
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 18432 5846 18460 10474
rect 19260 8566 19288 12786
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19904 10810 19932 10950
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19536 10062 19564 10678
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19628 9382 19656 10542
rect 20088 9586 20116 12582
rect 20272 10198 20300 18022
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18326 5536 18382 5545
rect 17899 5468 18195 5488
rect 18326 5471 18382 5480
rect 17955 5466 17979 5468
rect 18035 5466 18059 5468
rect 18115 5466 18139 5468
rect 17977 5414 17979 5466
rect 18041 5414 18053 5466
rect 18115 5414 18117 5466
rect 17955 5412 17979 5414
rect 18035 5412 18059 5414
rect 18115 5412 18139 5414
rect 17899 5392 18195 5412
rect 18340 5370 18368 5471
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 17899 4380 18195 4400
rect 17955 4378 17979 4380
rect 18035 4378 18059 4380
rect 18115 4378 18139 4380
rect 17977 4326 17979 4378
rect 18041 4326 18053 4378
rect 18115 4326 18117 4378
rect 17955 4324 17979 4326
rect 18035 4324 18059 4326
rect 18115 4324 18139 4326
rect 17899 4304 18195 4324
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 17899 3292 18195 3312
rect 17955 3290 17979 3292
rect 18035 3290 18059 3292
rect 18115 3290 18139 3292
rect 17977 3238 17979 3290
rect 18041 3238 18053 3290
rect 18115 3238 18117 3290
rect 17955 3236 17979 3238
rect 18035 3236 18059 3238
rect 18115 3236 18139 3238
rect 17899 3216 18195 3236
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 17899 2204 18195 2224
rect 17955 2202 17979 2204
rect 18035 2202 18059 2204
rect 18115 2202 18139 2204
rect 17977 2150 17979 2202
rect 18041 2150 18053 2202
rect 18115 2150 18117 2202
rect 17955 2148 17979 2150
rect 18035 2148 18059 2150
rect 18115 2148 18139 2150
rect 17899 2128 18195 2148
rect 19168 800 19196 4082
rect 570 0 626 800
rect 6642 0 6698 800
rect 12898 0 12954 800
rect 19154 0 19210 800
<< via2 >>
rect 2778 19080 2834 19136
rect 7733 22330 7789 22332
rect 7813 22330 7869 22332
rect 7893 22330 7949 22332
rect 7973 22330 8029 22332
rect 7733 22278 7759 22330
rect 7759 22278 7789 22330
rect 7813 22278 7823 22330
rect 7823 22278 7869 22330
rect 7893 22278 7939 22330
rect 7939 22278 7949 22330
rect 7973 22278 8003 22330
rect 8003 22278 8029 22330
rect 7733 22276 7789 22278
rect 7813 22276 7869 22278
rect 7893 22276 7949 22278
rect 7973 22276 8029 22278
rect 4344 21786 4400 21788
rect 4424 21786 4480 21788
rect 4504 21786 4560 21788
rect 4584 21786 4640 21788
rect 4344 21734 4370 21786
rect 4370 21734 4400 21786
rect 4424 21734 4434 21786
rect 4434 21734 4480 21786
rect 4504 21734 4550 21786
rect 4550 21734 4560 21786
rect 4584 21734 4614 21786
rect 4614 21734 4640 21786
rect 4344 21732 4400 21734
rect 4424 21732 4480 21734
rect 4504 21732 4560 21734
rect 4584 21732 4640 21734
rect 4344 20698 4400 20700
rect 4424 20698 4480 20700
rect 4504 20698 4560 20700
rect 4584 20698 4640 20700
rect 4344 20646 4370 20698
rect 4370 20646 4400 20698
rect 4424 20646 4434 20698
rect 4434 20646 4480 20698
rect 4504 20646 4550 20698
rect 4550 20646 4560 20698
rect 4584 20646 4614 20698
rect 4614 20646 4640 20698
rect 4344 20644 4400 20646
rect 4424 20644 4480 20646
rect 4504 20644 4560 20646
rect 4584 20644 4640 20646
rect 4344 19610 4400 19612
rect 4424 19610 4480 19612
rect 4504 19610 4560 19612
rect 4584 19610 4640 19612
rect 4344 19558 4370 19610
rect 4370 19558 4400 19610
rect 4424 19558 4434 19610
rect 4434 19558 4480 19610
rect 4504 19558 4550 19610
rect 4550 19558 4560 19610
rect 4584 19558 4614 19610
rect 4614 19558 4640 19610
rect 4344 19556 4400 19558
rect 4424 19556 4480 19558
rect 4504 19556 4560 19558
rect 4584 19556 4640 19558
rect 4344 18522 4400 18524
rect 4424 18522 4480 18524
rect 4504 18522 4560 18524
rect 4584 18522 4640 18524
rect 4344 18470 4370 18522
rect 4370 18470 4400 18522
rect 4424 18470 4434 18522
rect 4434 18470 4480 18522
rect 4504 18470 4550 18522
rect 4550 18470 4560 18522
rect 4584 18470 4614 18522
rect 4614 18470 4640 18522
rect 4344 18468 4400 18470
rect 4424 18468 4480 18470
rect 4504 18468 4560 18470
rect 4584 18468 4640 18470
rect 4344 17434 4400 17436
rect 4424 17434 4480 17436
rect 4504 17434 4560 17436
rect 4584 17434 4640 17436
rect 4344 17382 4370 17434
rect 4370 17382 4400 17434
rect 4424 17382 4434 17434
rect 4434 17382 4480 17434
rect 4504 17382 4550 17434
rect 4550 17382 4560 17434
rect 4584 17382 4614 17434
rect 4614 17382 4640 17434
rect 4344 17380 4400 17382
rect 4424 17380 4480 17382
rect 4504 17380 4560 17382
rect 4584 17380 4640 17382
rect 4344 16346 4400 16348
rect 4424 16346 4480 16348
rect 4504 16346 4560 16348
rect 4584 16346 4640 16348
rect 4344 16294 4370 16346
rect 4370 16294 4400 16346
rect 4424 16294 4434 16346
rect 4434 16294 4480 16346
rect 4504 16294 4550 16346
rect 4550 16294 4560 16346
rect 4584 16294 4614 16346
rect 4614 16294 4640 16346
rect 4344 16292 4400 16294
rect 4424 16292 4480 16294
rect 4504 16292 4560 16294
rect 4584 16292 4640 16294
rect 4344 15258 4400 15260
rect 4424 15258 4480 15260
rect 4504 15258 4560 15260
rect 4584 15258 4640 15260
rect 4344 15206 4370 15258
rect 4370 15206 4400 15258
rect 4424 15206 4434 15258
rect 4434 15206 4480 15258
rect 4504 15206 4550 15258
rect 4550 15206 4560 15258
rect 4584 15206 4614 15258
rect 4614 15206 4640 15258
rect 4344 15204 4400 15206
rect 4424 15204 4480 15206
rect 4504 15204 4560 15206
rect 4584 15204 4640 15206
rect 4344 14170 4400 14172
rect 4424 14170 4480 14172
rect 4504 14170 4560 14172
rect 4584 14170 4640 14172
rect 4344 14118 4370 14170
rect 4370 14118 4400 14170
rect 4424 14118 4434 14170
rect 4434 14118 4480 14170
rect 4504 14118 4550 14170
rect 4550 14118 4560 14170
rect 4584 14118 4614 14170
rect 4614 14118 4640 14170
rect 4344 14116 4400 14118
rect 4424 14116 4480 14118
rect 4504 14116 4560 14118
rect 4584 14116 4640 14118
rect 4344 13082 4400 13084
rect 4424 13082 4480 13084
rect 4504 13082 4560 13084
rect 4584 13082 4640 13084
rect 4344 13030 4370 13082
rect 4370 13030 4400 13082
rect 4424 13030 4434 13082
rect 4434 13030 4480 13082
rect 4504 13030 4550 13082
rect 4550 13030 4560 13082
rect 4584 13030 4614 13082
rect 4614 13030 4640 13082
rect 4344 13028 4400 13030
rect 4424 13028 4480 13030
rect 4504 13028 4560 13030
rect 4584 13028 4640 13030
rect 4344 11994 4400 11996
rect 4424 11994 4480 11996
rect 4504 11994 4560 11996
rect 4584 11994 4640 11996
rect 4344 11942 4370 11994
rect 4370 11942 4400 11994
rect 4424 11942 4434 11994
rect 4434 11942 4480 11994
rect 4504 11942 4550 11994
rect 4550 11942 4560 11994
rect 4584 11942 4614 11994
rect 4614 11942 4640 11994
rect 4344 11940 4400 11942
rect 4424 11940 4480 11942
rect 4504 11940 4560 11942
rect 4584 11940 4640 11942
rect 4344 10906 4400 10908
rect 4424 10906 4480 10908
rect 4504 10906 4560 10908
rect 4584 10906 4640 10908
rect 4344 10854 4370 10906
rect 4370 10854 4400 10906
rect 4424 10854 4434 10906
rect 4434 10854 4480 10906
rect 4504 10854 4550 10906
rect 4550 10854 4560 10906
rect 4584 10854 4614 10906
rect 4614 10854 4640 10906
rect 4344 10852 4400 10854
rect 4424 10852 4480 10854
rect 4504 10852 4560 10854
rect 4584 10852 4640 10854
rect 4066 9832 4122 9888
rect 4344 9818 4400 9820
rect 4424 9818 4480 9820
rect 4504 9818 4560 9820
rect 4584 9818 4640 9820
rect 4344 9766 4370 9818
rect 4370 9766 4400 9818
rect 4424 9766 4434 9818
rect 4434 9766 4480 9818
rect 4504 9766 4550 9818
rect 4550 9766 4560 9818
rect 4584 9766 4614 9818
rect 4614 9766 4640 9818
rect 4344 9764 4400 9766
rect 4424 9764 4480 9766
rect 4504 9764 4560 9766
rect 4584 9764 4640 9766
rect 4344 8730 4400 8732
rect 4424 8730 4480 8732
rect 4504 8730 4560 8732
rect 4584 8730 4640 8732
rect 4344 8678 4370 8730
rect 4370 8678 4400 8730
rect 4424 8678 4434 8730
rect 4434 8678 4480 8730
rect 4504 8678 4550 8730
rect 4550 8678 4560 8730
rect 4584 8678 4614 8730
rect 4614 8678 4640 8730
rect 4344 8676 4400 8678
rect 4424 8676 4480 8678
rect 4504 8676 4560 8678
rect 4584 8676 4640 8678
rect 4802 9696 4858 9752
rect 4344 7642 4400 7644
rect 4424 7642 4480 7644
rect 4504 7642 4560 7644
rect 4584 7642 4640 7644
rect 4344 7590 4370 7642
rect 4370 7590 4400 7642
rect 4424 7590 4434 7642
rect 4434 7590 4480 7642
rect 4504 7590 4550 7642
rect 4550 7590 4560 7642
rect 4584 7590 4614 7642
rect 4614 7590 4640 7642
rect 4344 7588 4400 7590
rect 4424 7588 4480 7590
rect 4504 7588 4560 7590
rect 4584 7588 4640 7590
rect 4344 6554 4400 6556
rect 4424 6554 4480 6556
rect 4504 6554 4560 6556
rect 4584 6554 4640 6556
rect 4344 6502 4370 6554
rect 4370 6502 4400 6554
rect 4424 6502 4434 6554
rect 4434 6502 4480 6554
rect 4504 6502 4550 6554
rect 4550 6502 4560 6554
rect 4584 6502 4614 6554
rect 4614 6502 4640 6554
rect 4344 6500 4400 6502
rect 4424 6500 4480 6502
rect 4504 6500 4560 6502
rect 4584 6500 4640 6502
rect 4344 5466 4400 5468
rect 4424 5466 4480 5468
rect 4504 5466 4560 5468
rect 4584 5466 4640 5468
rect 4344 5414 4370 5466
rect 4370 5414 4400 5466
rect 4424 5414 4434 5466
rect 4434 5414 4480 5466
rect 4504 5414 4550 5466
rect 4550 5414 4560 5466
rect 4584 5414 4614 5466
rect 4614 5414 4640 5466
rect 4344 5412 4400 5414
rect 4424 5412 4480 5414
rect 4504 5412 4560 5414
rect 4584 5412 4640 5414
rect 4344 4378 4400 4380
rect 4424 4378 4480 4380
rect 4504 4378 4560 4380
rect 4584 4378 4640 4380
rect 4344 4326 4370 4378
rect 4370 4326 4400 4378
rect 4424 4326 4434 4378
rect 4434 4326 4480 4378
rect 4504 4326 4550 4378
rect 4550 4326 4560 4378
rect 4584 4326 4614 4378
rect 4614 4326 4640 4378
rect 4344 4324 4400 4326
rect 4424 4324 4480 4326
rect 4504 4324 4560 4326
rect 4584 4324 4640 4326
rect 4344 3290 4400 3292
rect 4424 3290 4480 3292
rect 4504 3290 4560 3292
rect 4584 3290 4640 3292
rect 4344 3238 4370 3290
rect 4370 3238 4400 3290
rect 4424 3238 4434 3290
rect 4434 3238 4480 3290
rect 4504 3238 4550 3290
rect 4550 3238 4560 3290
rect 4584 3238 4614 3290
rect 4614 3238 4640 3290
rect 4344 3236 4400 3238
rect 4424 3236 4480 3238
rect 4504 3236 4560 3238
rect 4584 3236 4640 3238
rect 5354 9696 5410 9752
rect 7733 21242 7789 21244
rect 7813 21242 7869 21244
rect 7893 21242 7949 21244
rect 7973 21242 8029 21244
rect 7733 21190 7759 21242
rect 7759 21190 7789 21242
rect 7813 21190 7823 21242
rect 7823 21190 7869 21242
rect 7893 21190 7939 21242
rect 7939 21190 7949 21242
rect 7973 21190 8003 21242
rect 8003 21190 8029 21242
rect 7733 21188 7789 21190
rect 7813 21188 7869 21190
rect 7893 21188 7949 21190
rect 7973 21188 8029 21190
rect 7733 20154 7789 20156
rect 7813 20154 7869 20156
rect 7893 20154 7949 20156
rect 7973 20154 8029 20156
rect 7733 20102 7759 20154
rect 7759 20102 7789 20154
rect 7813 20102 7823 20154
rect 7823 20102 7869 20154
rect 7893 20102 7939 20154
rect 7939 20102 7949 20154
rect 7973 20102 8003 20154
rect 8003 20102 8029 20154
rect 7733 20100 7789 20102
rect 7813 20100 7869 20102
rect 7893 20100 7949 20102
rect 7973 20100 8029 20102
rect 7733 19066 7789 19068
rect 7813 19066 7869 19068
rect 7893 19066 7949 19068
rect 7973 19066 8029 19068
rect 7733 19014 7759 19066
rect 7759 19014 7789 19066
rect 7813 19014 7823 19066
rect 7823 19014 7869 19066
rect 7893 19014 7939 19066
rect 7939 19014 7949 19066
rect 7973 19014 8003 19066
rect 8003 19014 8029 19066
rect 7733 19012 7789 19014
rect 7813 19012 7869 19014
rect 7893 19012 7949 19014
rect 7973 19012 8029 19014
rect 4344 2202 4400 2204
rect 4424 2202 4480 2204
rect 4504 2202 4560 2204
rect 4584 2202 4640 2204
rect 4344 2150 4370 2202
rect 4370 2150 4400 2202
rect 4424 2150 4434 2202
rect 4434 2150 4480 2202
rect 4504 2150 4550 2202
rect 4550 2150 4560 2202
rect 4584 2150 4614 2202
rect 4614 2150 4640 2202
rect 4344 2148 4400 2150
rect 4424 2148 4480 2150
rect 4504 2148 4560 2150
rect 4584 2148 4640 2150
rect 7733 17978 7789 17980
rect 7813 17978 7869 17980
rect 7893 17978 7949 17980
rect 7973 17978 8029 17980
rect 7733 17926 7759 17978
rect 7759 17926 7789 17978
rect 7813 17926 7823 17978
rect 7823 17926 7869 17978
rect 7893 17926 7939 17978
rect 7939 17926 7949 17978
rect 7973 17926 8003 17978
rect 8003 17926 8029 17978
rect 7733 17924 7789 17926
rect 7813 17924 7869 17926
rect 7893 17924 7949 17926
rect 7973 17924 8029 17926
rect 7733 16890 7789 16892
rect 7813 16890 7869 16892
rect 7893 16890 7949 16892
rect 7973 16890 8029 16892
rect 7733 16838 7759 16890
rect 7759 16838 7789 16890
rect 7813 16838 7823 16890
rect 7823 16838 7869 16890
rect 7893 16838 7939 16890
rect 7939 16838 7949 16890
rect 7973 16838 8003 16890
rect 8003 16838 8029 16890
rect 7733 16836 7789 16838
rect 7813 16836 7869 16838
rect 7893 16836 7949 16838
rect 7973 16836 8029 16838
rect 7733 15802 7789 15804
rect 7813 15802 7869 15804
rect 7893 15802 7949 15804
rect 7973 15802 8029 15804
rect 7733 15750 7759 15802
rect 7759 15750 7789 15802
rect 7813 15750 7823 15802
rect 7823 15750 7869 15802
rect 7893 15750 7939 15802
rect 7939 15750 7949 15802
rect 7973 15750 8003 15802
rect 8003 15750 8029 15802
rect 7733 15748 7789 15750
rect 7813 15748 7869 15750
rect 7893 15748 7949 15750
rect 7973 15748 8029 15750
rect 7733 14714 7789 14716
rect 7813 14714 7869 14716
rect 7893 14714 7949 14716
rect 7973 14714 8029 14716
rect 7733 14662 7759 14714
rect 7759 14662 7789 14714
rect 7813 14662 7823 14714
rect 7823 14662 7869 14714
rect 7893 14662 7939 14714
rect 7939 14662 7949 14714
rect 7973 14662 8003 14714
rect 8003 14662 8029 14714
rect 7733 14660 7789 14662
rect 7813 14660 7869 14662
rect 7893 14660 7949 14662
rect 7973 14660 8029 14662
rect 7733 13626 7789 13628
rect 7813 13626 7869 13628
rect 7893 13626 7949 13628
rect 7973 13626 8029 13628
rect 7733 13574 7759 13626
rect 7759 13574 7789 13626
rect 7813 13574 7823 13626
rect 7823 13574 7869 13626
rect 7893 13574 7939 13626
rect 7939 13574 7949 13626
rect 7973 13574 8003 13626
rect 8003 13574 8029 13626
rect 7733 13572 7789 13574
rect 7813 13572 7869 13574
rect 7893 13572 7949 13574
rect 7973 13572 8029 13574
rect 7733 12538 7789 12540
rect 7813 12538 7869 12540
rect 7893 12538 7949 12540
rect 7973 12538 8029 12540
rect 7733 12486 7759 12538
rect 7759 12486 7789 12538
rect 7813 12486 7823 12538
rect 7823 12486 7869 12538
rect 7893 12486 7939 12538
rect 7939 12486 7949 12538
rect 7973 12486 8003 12538
rect 8003 12486 8029 12538
rect 7733 12484 7789 12486
rect 7813 12484 7869 12486
rect 7893 12484 7949 12486
rect 7973 12484 8029 12486
rect 7733 11450 7789 11452
rect 7813 11450 7869 11452
rect 7893 11450 7949 11452
rect 7973 11450 8029 11452
rect 7733 11398 7759 11450
rect 7759 11398 7789 11450
rect 7813 11398 7823 11450
rect 7823 11398 7869 11450
rect 7893 11398 7939 11450
rect 7939 11398 7949 11450
rect 7973 11398 8003 11450
rect 8003 11398 8029 11450
rect 7733 11396 7789 11398
rect 7813 11396 7869 11398
rect 7893 11396 7949 11398
rect 7973 11396 8029 11398
rect 7733 10362 7789 10364
rect 7813 10362 7869 10364
rect 7893 10362 7949 10364
rect 7973 10362 8029 10364
rect 7733 10310 7759 10362
rect 7759 10310 7789 10362
rect 7813 10310 7823 10362
rect 7823 10310 7869 10362
rect 7893 10310 7939 10362
rect 7939 10310 7949 10362
rect 7973 10310 8003 10362
rect 8003 10310 8029 10362
rect 7733 10308 7789 10310
rect 7813 10308 7869 10310
rect 7893 10308 7949 10310
rect 7973 10308 8029 10310
rect 7733 9274 7789 9276
rect 7813 9274 7869 9276
rect 7893 9274 7949 9276
rect 7973 9274 8029 9276
rect 7733 9222 7759 9274
rect 7759 9222 7789 9274
rect 7813 9222 7823 9274
rect 7823 9222 7869 9274
rect 7893 9222 7939 9274
rect 7939 9222 7949 9274
rect 7973 9222 8003 9274
rect 8003 9222 8029 9274
rect 7733 9220 7789 9222
rect 7813 9220 7869 9222
rect 7893 9220 7949 9222
rect 7973 9220 8029 9222
rect 7733 8186 7789 8188
rect 7813 8186 7869 8188
rect 7893 8186 7949 8188
rect 7973 8186 8029 8188
rect 7733 8134 7759 8186
rect 7759 8134 7789 8186
rect 7813 8134 7823 8186
rect 7823 8134 7869 8186
rect 7893 8134 7939 8186
rect 7939 8134 7949 8186
rect 7973 8134 8003 8186
rect 8003 8134 8029 8186
rect 7733 8132 7789 8134
rect 7813 8132 7869 8134
rect 7893 8132 7949 8134
rect 7973 8132 8029 8134
rect 7733 7098 7789 7100
rect 7813 7098 7869 7100
rect 7893 7098 7949 7100
rect 7973 7098 8029 7100
rect 7733 7046 7759 7098
rect 7759 7046 7789 7098
rect 7813 7046 7823 7098
rect 7823 7046 7869 7098
rect 7893 7046 7939 7098
rect 7939 7046 7949 7098
rect 7973 7046 8003 7098
rect 8003 7046 8029 7098
rect 7733 7044 7789 7046
rect 7813 7044 7869 7046
rect 7893 7044 7949 7046
rect 7973 7044 8029 7046
rect 7733 6010 7789 6012
rect 7813 6010 7869 6012
rect 7893 6010 7949 6012
rect 7973 6010 8029 6012
rect 7733 5958 7759 6010
rect 7759 5958 7789 6010
rect 7813 5958 7823 6010
rect 7823 5958 7869 6010
rect 7893 5958 7939 6010
rect 7939 5958 7949 6010
rect 7973 5958 8003 6010
rect 8003 5958 8029 6010
rect 7733 5956 7789 5958
rect 7813 5956 7869 5958
rect 7893 5956 7949 5958
rect 7973 5956 8029 5958
rect 7733 4922 7789 4924
rect 7813 4922 7869 4924
rect 7893 4922 7949 4924
rect 7973 4922 8029 4924
rect 7733 4870 7759 4922
rect 7759 4870 7789 4922
rect 7813 4870 7823 4922
rect 7823 4870 7869 4922
rect 7893 4870 7939 4922
rect 7939 4870 7949 4922
rect 7973 4870 8003 4922
rect 8003 4870 8029 4922
rect 7733 4868 7789 4870
rect 7813 4868 7869 4870
rect 7893 4868 7949 4870
rect 7973 4868 8029 4870
rect 7733 3834 7789 3836
rect 7813 3834 7869 3836
rect 7893 3834 7949 3836
rect 7973 3834 8029 3836
rect 7733 3782 7759 3834
rect 7759 3782 7789 3834
rect 7813 3782 7823 3834
rect 7823 3782 7869 3834
rect 7893 3782 7939 3834
rect 7939 3782 7949 3834
rect 7973 3782 8003 3834
rect 8003 3782 8029 3834
rect 7733 3780 7789 3782
rect 7813 3780 7869 3782
rect 7893 3780 7949 3782
rect 7973 3780 8029 3782
rect 7733 2746 7789 2748
rect 7813 2746 7869 2748
rect 7893 2746 7949 2748
rect 7973 2746 8029 2748
rect 7733 2694 7759 2746
rect 7759 2694 7789 2746
rect 7813 2694 7823 2746
rect 7823 2694 7869 2746
rect 7893 2694 7939 2746
rect 7939 2694 7949 2746
rect 7973 2694 8003 2746
rect 8003 2694 8029 2746
rect 7733 2692 7789 2694
rect 7813 2692 7869 2694
rect 7893 2692 7949 2694
rect 7973 2692 8029 2694
rect 14510 22330 14566 22332
rect 14590 22330 14646 22332
rect 14670 22330 14726 22332
rect 14750 22330 14806 22332
rect 14510 22278 14536 22330
rect 14536 22278 14566 22330
rect 14590 22278 14600 22330
rect 14600 22278 14646 22330
rect 14670 22278 14716 22330
rect 14716 22278 14726 22330
rect 14750 22278 14780 22330
rect 14780 22278 14806 22330
rect 14510 22276 14566 22278
rect 14590 22276 14646 22278
rect 14670 22276 14726 22278
rect 14750 22276 14806 22278
rect 11122 21786 11178 21788
rect 11202 21786 11258 21788
rect 11282 21786 11338 21788
rect 11362 21786 11418 21788
rect 11122 21734 11148 21786
rect 11148 21734 11178 21786
rect 11202 21734 11212 21786
rect 11212 21734 11258 21786
rect 11282 21734 11328 21786
rect 11328 21734 11338 21786
rect 11362 21734 11392 21786
rect 11392 21734 11418 21786
rect 11122 21732 11178 21734
rect 11202 21732 11258 21734
rect 11282 21732 11338 21734
rect 11362 21732 11418 21734
rect 11122 20698 11178 20700
rect 11202 20698 11258 20700
rect 11282 20698 11338 20700
rect 11362 20698 11418 20700
rect 11122 20646 11148 20698
rect 11148 20646 11178 20698
rect 11202 20646 11212 20698
rect 11212 20646 11258 20698
rect 11282 20646 11328 20698
rect 11328 20646 11338 20698
rect 11362 20646 11392 20698
rect 11392 20646 11418 20698
rect 11122 20644 11178 20646
rect 11202 20644 11258 20646
rect 11282 20644 11338 20646
rect 11362 20644 11418 20646
rect 11122 19610 11178 19612
rect 11202 19610 11258 19612
rect 11282 19610 11338 19612
rect 11362 19610 11418 19612
rect 11122 19558 11148 19610
rect 11148 19558 11178 19610
rect 11202 19558 11212 19610
rect 11212 19558 11258 19610
rect 11282 19558 11328 19610
rect 11328 19558 11338 19610
rect 11362 19558 11392 19610
rect 11392 19558 11418 19610
rect 11122 19556 11178 19558
rect 11202 19556 11258 19558
rect 11282 19556 11338 19558
rect 11362 19556 11418 19558
rect 11122 18522 11178 18524
rect 11202 18522 11258 18524
rect 11282 18522 11338 18524
rect 11362 18522 11418 18524
rect 11122 18470 11148 18522
rect 11148 18470 11178 18522
rect 11202 18470 11212 18522
rect 11212 18470 11258 18522
rect 11282 18470 11328 18522
rect 11328 18470 11338 18522
rect 11362 18470 11392 18522
rect 11392 18470 11418 18522
rect 11122 18468 11178 18470
rect 11202 18468 11258 18470
rect 11282 18468 11338 18470
rect 11362 18468 11418 18470
rect 11122 17434 11178 17436
rect 11202 17434 11258 17436
rect 11282 17434 11338 17436
rect 11362 17434 11418 17436
rect 11122 17382 11148 17434
rect 11148 17382 11178 17434
rect 11202 17382 11212 17434
rect 11212 17382 11258 17434
rect 11282 17382 11328 17434
rect 11328 17382 11338 17434
rect 11362 17382 11392 17434
rect 11392 17382 11418 17434
rect 11122 17380 11178 17382
rect 11202 17380 11258 17382
rect 11282 17380 11338 17382
rect 11362 17380 11418 17382
rect 11122 16346 11178 16348
rect 11202 16346 11258 16348
rect 11282 16346 11338 16348
rect 11362 16346 11418 16348
rect 11122 16294 11148 16346
rect 11148 16294 11178 16346
rect 11202 16294 11212 16346
rect 11212 16294 11258 16346
rect 11282 16294 11328 16346
rect 11328 16294 11338 16346
rect 11362 16294 11392 16346
rect 11392 16294 11418 16346
rect 11122 16292 11178 16294
rect 11202 16292 11258 16294
rect 11282 16292 11338 16294
rect 11362 16292 11418 16294
rect 11122 15258 11178 15260
rect 11202 15258 11258 15260
rect 11282 15258 11338 15260
rect 11362 15258 11418 15260
rect 11122 15206 11148 15258
rect 11148 15206 11178 15258
rect 11202 15206 11212 15258
rect 11212 15206 11258 15258
rect 11282 15206 11328 15258
rect 11328 15206 11338 15258
rect 11362 15206 11392 15258
rect 11392 15206 11418 15258
rect 11122 15204 11178 15206
rect 11202 15204 11258 15206
rect 11282 15204 11338 15206
rect 11362 15204 11418 15206
rect 11122 14170 11178 14172
rect 11202 14170 11258 14172
rect 11282 14170 11338 14172
rect 11362 14170 11418 14172
rect 11122 14118 11148 14170
rect 11148 14118 11178 14170
rect 11202 14118 11212 14170
rect 11212 14118 11258 14170
rect 11282 14118 11328 14170
rect 11328 14118 11338 14170
rect 11362 14118 11392 14170
rect 11392 14118 11418 14170
rect 11122 14116 11178 14118
rect 11202 14116 11258 14118
rect 11282 14116 11338 14118
rect 11362 14116 11418 14118
rect 11122 13082 11178 13084
rect 11202 13082 11258 13084
rect 11282 13082 11338 13084
rect 11362 13082 11418 13084
rect 11122 13030 11148 13082
rect 11148 13030 11178 13082
rect 11202 13030 11212 13082
rect 11212 13030 11258 13082
rect 11282 13030 11328 13082
rect 11328 13030 11338 13082
rect 11362 13030 11392 13082
rect 11392 13030 11418 13082
rect 11122 13028 11178 13030
rect 11202 13028 11258 13030
rect 11282 13028 11338 13030
rect 11362 13028 11418 13030
rect 11122 11994 11178 11996
rect 11202 11994 11258 11996
rect 11282 11994 11338 11996
rect 11362 11994 11418 11996
rect 11122 11942 11148 11994
rect 11148 11942 11178 11994
rect 11202 11942 11212 11994
rect 11212 11942 11258 11994
rect 11282 11942 11328 11994
rect 11328 11942 11338 11994
rect 11362 11942 11392 11994
rect 11392 11942 11418 11994
rect 11122 11940 11178 11942
rect 11202 11940 11258 11942
rect 11282 11940 11338 11942
rect 11362 11940 11418 11942
rect 11122 10906 11178 10908
rect 11202 10906 11258 10908
rect 11282 10906 11338 10908
rect 11362 10906 11418 10908
rect 11122 10854 11148 10906
rect 11148 10854 11178 10906
rect 11202 10854 11212 10906
rect 11212 10854 11258 10906
rect 11282 10854 11328 10906
rect 11328 10854 11338 10906
rect 11362 10854 11392 10906
rect 11392 10854 11418 10906
rect 11122 10852 11178 10854
rect 11202 10852 11258 10854
rect 11282 10852 11338 10854
rect 11362 10852 11418 10854
rect 11122 9818 11178 9820
rect 11202 9818 11258 9820
rect 11282 9818 11338 9820
rect 11362 9818 11418 9820
rect 11122 9766 11148 9818
rect 11148 9766 11178 9818
rect 11202 9766 11212 9818
rect 11212 9766 11258 9818
rect 11282 9766 11328 9818
rect 11328 9766 11338 9818
rect 11362 9766 11392 9818
rect 11392 9766 11418 9818
rect 11122 9764 11178 9766
rect 11202 9764 11258 9766
rect 11282 9764 11338 9766
rect 11362 9764 11418 9766
rect 11122 8730 11178 8732
rect 11202 8730 11258 8732
rect 11282 8730 11338 8732
rect 11362 8730 11418 8732
rect 11122 8678 11148 8730
rect 11148 8678 11178 8730
rect 11202 8678 11212 8730
rect 11212 8678 11258 8730
rect 11282 8678 11328 8730
rect 11328 8678 11338 8730
rect 11362 8678 11392 8730
rect 11392 8678 11418 8730
rect 11122 8676 11178 8678
rect 11202 8676 11258 8678
rect 11282 8676 11338 8678
rect 11362 8676 11418 8678
rect 11122 7642 11178 7644
rect 11202 7642 11258 7644
rect 11282 7642 11338 7644
rect 11362 7642 11418 7644
rect 11122 7590 11148 7642
rect 11148 7590 11178 7642
rect 11202 7590 11212 7642
rect 11212 7590 11258 7642
rect 11282 7590 11328 7642
rect 11328 7590 11338 7642
rect 11362 7590 11392 7642
rect 11392 7590 11418 7642
rect 11122 7588 11178 7590
rect 11202 7588 11258 7590
rect 11282 7588 11338 7590
rect 11362 7588 11418 7590
rect 11122 6554 11178 6556
rect 11202 6554 11258 6556
rect 11282 6554 11338 6556
rect 11362 6554 11418 6556
rect 11122 6502 11148 6554
rect 11148 6502 11178 6554
rect 11202 6502 11212 6554
rect 11212 6502 11258 6554
rect 11282 6502 11328 6554
rect 11328 6502 11338 6554
rect 11362 6502 11392 6554
rect 11392 6502 11418 6554
rect 11122 6500 11178 6502
rect 11202 6500 11258 6502
rect 11282 6500 11338 6502
rect 11362 6500 11418 6502
rect 11122 5466 11178 5468
rect 11202 5466 11258 5468
rect 11282 5466 11338 5468
rect 11362 5466 11418 5468
rect 11122 5414 11148 5466
rect 11148 5414 11178 5466
rect 11202 5414 11212 5466
rect 11212 5414 11258 5466
rect 11282 5414 11328 5466
rect 11328 5414 11338 5466
rect 11362 5414 11392 5466
rect 11392 5414 11418 5466
rect 11122 5412 11178 5414
rect 11202 5412 11258 5414
rect 11282 5412 11338 5414
rect 11362 5412 11418 5414
rect 11122 4378 11178 4380
rect 11202 4378 11258 4380
rect 11282 4378 11338 4380
rect 11362 4378 11418 4380
rect 11122 4326 11148 4378
rect 11148 4326 11178 4378
rect 11202 4326 11212 4378
rect 11212 4326 11258 4378
rect 11282 4326 11328 4378
rect 11328 4326 11338 4378
rect 11362 4326 11392 4378
rect 11392 4326 11418 4378
rect 11122 4324 11178 4326
rect 11202 4324 11258 4326
rect 11282 4324 11338 4326
rect 11362 4324 11418 4326
rect 11122 3290 11178 3292
rect 11202 3290 11258 3292
rect 11282 3290 11338 3292
rect 11362 3290 11418 3292
rect 11122 3238 11148 3290
rect 11148 3238 11178 3290
rect 11202 3238 11212 3290
rect 11212 3238 11258 3290
rect 11282 3238 11328 3290
rect 11328 3238 11338 3290
rect 11362 3238 11392 3290
rect 11392 3238 11418 3290
rect 11122 3236 11178 3238
rect 11202 3236 11258 3238
rect 11282 3236 11338 3238
rect 11362 3236 11418 3238
rect 12622 9594 12678 9650
rect 14510 21242 14566 21244
rect 14590 21242 14646 21244
rect 14670 21242 14726 21244
rect 14750 21242 14806 21244
rect 14510 21190 14536 21242
rect 14536 21190 14566 21242
rect 14590 21190 14600 21242
rect 14600 21190 14646 21242
rect 14670 21190 14716 21242
rect 14716 21190 14726 21242
rect 14750 21190 14780 21242
rect 14780 21190 14806 21242
rect 14510 21188 14566 21190
rect 14590 21188 14646 21190
rect 14670 21188 14726 21190
rect 14750 21188 14806 21190
rect 14510 20154 14566 20156
rect 14590 20154 14646 20156
rect 14670 20154 14726 20156
rect 14750 20154 14806 20156
rect 14510 20102 14536 20154
rect 14536 20102 14566 20154
rect 14590 20102 14600 20154
rect 14600 20102 14646 20154
rect 14670 20102 14716 20154
rect 14716 20102 14726 20154
rect 14750 20102 14780 20154
rect 14780 20102 14806 20154
rect 14510 20100 14566 20102
rect 14590 20100 14646 20102
rect 14670 20100 14726 20102
rect 14750 20100 14806 20102
rect 14510 19066 14566 19068
rect 14590 19066 14646 19068
rect 14670 19066 14726 19068
rect 14750 19066 14806 19068
rect 14510 19014 14536 19066
rect 14536 19014 14566 19066
rect 14590 19014 14600 19066
rect 14600 19014 14646 19066
rect 14670 19014 14716 19066
rect 14716 19014 14726 19066
rect 14750 19014 14780 19066
rect 14780 19014 14806 19066
rect 14510 19012 14566 19014
rect 14590 19012 14646 19014
rect 14670 19012 14726 19014
rect 14750 19012 14806 19014
rect 14510 17978 14566 17980
rect 14590 17978 14646 17980
rect 14670 17978 14726 17980
rect 14750 17978 14806 17980
rect 14510 17926 14536 17978
rect 14536 17926 14566 17978
rect 14590 17926 14600 17978
rect 14600 17926 14646 17978
rect 14670 17926 14716 17978
rect 14716 17926 14726 17978
rect 14750 17926 14780 17978
rect 14780 17926 14806 17978
rect 14510 17924 14566 17926
rect 14590 17924 14646 17926
rect 14670 17924 14726 17926
rect 14750 17924 14806 17926
rect 13266 9696 13322 9752
rect 12990 9560 13046 9616
rect 12898 8492 12954 8528
rect 12898 8472 12900 8492
rect 12900 8472 12952 8492
rect 12952 8472 12954 8492
rect 11122 2202 11178 2204
rect 11202 2202 11258 2204
rect 11282 2202 11338 2204
rect 11362 2202 11418 2204
rect 11122 2150 11148 2202
rect 11148 2150 11178 2202
rect 11202 2150 11212 2202
rect 11212 2150 11258 2202
rect 11282 2150 11328 2202
rect 11328 2150 11338 2202
rect 11362 2150 11392 2202
rect 11392 2150 11418 2202
rect 11122 2148 11178 2150
rect 11202 2148 11258 2150
rect 11282 2148 11338 2150
rect 11362 2148 11418 2150
rect 14510 16890 14566 16892
rect 14590 16890 14646 16892
rect 14670 16890 14726 16892
rect 14750 16890 14806 16892
rect 14510 16838 14536 16890
rect 14536 16838 14566 16890
rect 14590 16838 14600 16890
rect 14600 16838 14646 16890
rect 14670 16838 14716 16890
rect 14716 16838 14726 16890
rect 14750 16838 14780 16890
rect 14780 16838 14806 16890
rect 14510 16836 14566 16838
rect 14590 16836 14646 16838
rect 14670 16836 14726 16838
rect 14750 16836 14806 16838
rect 14510 15802 14566 15804
rect 14590 15802 14646 15804
rect 14670 15802 14726 15804
rect 14750 15802 14806 15804
rect 14510 15750 14536 15802
rect 14536 15750 14566 15802
rect 14590 15750 14600 15802
rect 14600 15750 14646 15802
rect 14670 15750 14716 15802
rect 14716 15750 14726 15802
rect 14750 15750 14780 15802
rect 14780 15750 14806 15802
rect 14510 15748 14566 15750
rect 14590 15748 14646 15750
rect 14670 15748 14726 15750
rect 14750 15748 14806 15750
rect 14510 14714 14566 14716
rect 14590 14714 14646 14716
rect 14670 14714 14726 14716
rect 14750 14714 14806 14716
rect 14510 14662 14536 14714
rect 14536 14662 14566 14714
rect 14590 14662 14600 14714
rect 14600 14662 14646 14714
rect 14670 14662 14716 14714
rect 14716 14662 14726 14714
rect 14750 14662 14780 14714
rect 14780 14662 14806 14714
rect 14510 14660 14566 14662
rect 14590 14660 14646 14662
rect 14670 14660 14726 14662
rect 14750 14660 14806 14662
rect 14510 13626 14566 13628
rect 14590 13626 14646 13628
rect 14670 13626 14726 13628
rect 14750 13626 14806 13628
rect 14510 13574 14536 13626
rect 14536 13574 14566 13626
rect 14590 13574 14600 13626
rect 14600 13574 14646 13626
rect 14670 13574 14716 13626
rect 14716 13574 14726 13626
rect 14750 13574 14780 13626
rect 14780 13574 14806 13626
rect 14510 13572 14566 13574
rect 14590 13572 14646 13574
rect 14670 13572 14726 13574
rect 14750 13572 14806 13574
rect 14510 12538 14566 12540
rect 14590 12538 14646 12540
rect 14670 12538 14726 12540
rect 14750 12538 14806 12540
rect 14510 12486 14536 12538
rect 14536 12486 14566 12538
rect 14590 12486 14600 12538
rect 14600 12486 14646 12538
rect 14670 12486 14716 12538
rect 14716 12486 14726 12538
rect 14750 12486 14780 12538
rect 14780 12486 14806 12538
rect 14510 12484 14566 12486
rect 14590 12484 14646 12486
rect 14670 12484 14726 12486
rect 14750 12484 14806 12486
rect 14510 11450 14566 11452
rect 14590 11450 14646 11452
rect 14670 11450 14726 11452
rect 14750 11450 14806 11452
rect 14510 11398 14536 11450
rect 14536 11398 14566 11450
rect 14590 11398 14600 11450
rect 14600 11398 14646 11450
rect 14670 11398 14716 11450
rect 14716 11398 14726 11450
rect 14750 11398 14780 11450
rect 14780 11398 14806 11450
rect 14510 11396 14566 11398
rect 14590 11396 14646 11398
rect 14670 11396 14726 11398
rect 14750 11396 14806 11398
rect 14510 10362 14566 10364
rect 14590 10362 14646 10364
rect 14670 10362 14726 10364
rect 14750 10362 14806 10364
rect 14510 10310 14536 10362
rect 14536 10310 14566 10362
rect 14590 10310 14600 10362
rect 14600 10310 14646 10362
rect 14670 10310 14716 10362
rect 14716 10310 14726 10362
rect 14750 10310 14780 10362
rect 14780 10310 14806 10362
rect 14510 10308 14566 10310
rect 14590 10308 14646 10310
rect 14670 10308 14726 10310
rect 14750 10308 14806 10310
rect 14510 9274 14566 9276
rect 14590 9274 14646 9276
rect 14670 9274 14726 9276
rect 14750 9274 14806 9276
rect 14510 9222 14536 9274
rect 14536 9222 14566 9274
rect 14590 9222 14600 9274
rect 14600 9222 14646 9274
rect 14670 9222 14716 9274
rect 14716 9222 14726 9274
rect 14750 9222 14780 9274
rect 14780 9222 14806 9274
rect 14510 9220 14566 9222
rect 14590 9220 14646 9222
rect 14670 9220 14726 9222
rect 14750 9220 14806 9222
rect 17899 21786 17955 21788
rect 17979 21786 18035 21788
rect 18059 21786 18115 21788
rect 18139 21786 18195 21788
rect 17899 21734 17925 21786
rect 17925 21734 17955 21786
rect 17979 21734 17989 21786
rect 17989 21734 18035 21786
rect 18059 21734 18105 21786
rect 18105 21734 18115 21786
rect 18139 21734 18169 21786
rect 18169 21734 18195 21786
rect 17899 21732 17955 21734
rect 17979 21732 18035 21734
rect 18059 21732 18115 21734
rect 18139 21732 18195 21734
rect 14510 8186 14566 8188
rect 14590 8186 14646 8188
rect 14670 8186 14726 8188
rect 14750 8186 14806 8188
rect 14510 8134 14536 8186
rect 14536 8134 14566 8186
rect 14590 8134 14600 8186
rect 14600 8134 14646 8186
rect 14670 8134 14716 8186
rect 14716 8134 14726 8186
rect 14750 8134 14780 8186
rect 14780 8134 14806 8186
rect 14510 8132 14566 8134
rect 14590 8132 14646 8134
rect 14670 8132 14726 8134
rect 14750 8132 14806 8134
rect 14510 7098 14566 7100
rect 14590 7098 14646 7100
rect 14670 7098 14726 7100
rect 14750 7098 14806 7100
rect 14510 7046 14536 7098
rect 14536 7046 14566 7098
rect 14590 7046 14600 7098
rect 14600 7046 14646 7098
rect 14670 7046 14716 7098
rect 14716 7046 14726 7098
rect 14750 7046 14780 7098
rect 14780 7046 14806 7098
rect 14510 7044 14566 7046
rect 14590 7044 14646 7046
rect 14670 7044 14726 7046
rect 14750 7044 14806 7046
rect 14510 6010 14566 6012
rect 14590 6010 14646 6012
rect 14670 6010 14726 6012
rect 14750 6010 14806 6012
rect 14510 5958 14536 6010
rect 14536 5958 14566 6010
rect 14590 5958 14600 6010
rect 14600 5958 14646 6010
rect 14670 5958 14716 6010
rect 14716 5958 14726 6010
rect 14750 5958 14780 6010
rect 14780 5958 14806 6010
rect 14510 5956 14566 5958
rect 14590 5956 14646 5958
rect 14670 5956 14726 5958
rect 14750 5956 14806 5958
rect 14510 4922 14566 4924
rect 14590 4922 14646 4924
rect 14670 4922 14726 4924
rect 14750 4922 14806 4924
rect 14510 4870 14536 4922
rect 14536 4870 14566 4922
rect 14590 4870 14600 4922
rect 14600 4870 14646 4922
rect 14670 4870 14716 4922
rect 14716 4870 14726 4922
rect 14750 4870 14780 4922
rect 14780 4870 14806 4922
rect 14510 4868 14566 4870
rect 14590 4868 14646 4870
rect 14670 4868 14726 4870
rect 14750 4868 14806 4870
rect 14510 3834 14566 3836
rect 14590 3834 14646 3836
rect 14670 3834 14726 3836
rect 14750 3834 14806 3836
rect 14510 3782 14536 3834
rect 14536 3782 14566 3834
rect 14590 3782 14600 3834
rect 14600 3782 14646 3834
rect 14670 3782 14716 3834
rect 14716 3782 14726 3834
rect 14750 3782 14780 3834
rect 14780 3782 14806 3834
rect 14510 3780 14566 3782
rect 14590 3780 14646 3782
rect 14670 3780 14726 3782
rect 14750 3780 14806 3782
rect 15842 9560 15898 9616
rect 15750 8492 15806 8528
rect 15750 8472 15752 8492
rect 15752 8472 15804 8492
rect 15804 8472 15806 8492
rect 14510 2746 14566 2748
rect 14590 2746 14646 2748
rect 14670 2746 14726 2748
rect 14750 2746 14806 2748
rect 14510 2694 14536 2746
rect 14536 2694 14566 2746
rect 14590 2694 14600 2746
rect 14600 2694 14646 2746
rect 14670 2694 14716 2746
rect 14716 2694 14726 2746
rect 14750 2694 14780 2746
rect 14780 2694 14806 2746
rect 14510 2692 14566 2694
rect 14590 2692 14646 2694
rect 14670 2692 14726 2694
rect 14750 2692 14806 2694
rect 17899 20698 17955 20700
rect 17979 20698 18035 20700
rect 18059 20698 18115 20700
rect 18139 20698 18195 20700
rect 17899 20646 17925 20698
rect 17925 20646 17955 20698
rect 17979 20646 17989 20698
rect 17989 20646 18035 20698
rect 18059 20646 18105 20698
rect 18105 20646 18115 20698
rect 18139 20646 18169 20698
rect 18169 20646 18195 20698
rect 17899 20644 17955 20646
rect 17979 20644 18035 20646
rect 18059 20644 18115 20646
rect 18139 20644 18195 20646
rect 17899 19610 17955 19612
rect 17979 19610 18035 19612
rect 18059 19610 18115 19612
rect 18139 19610 18195 19612
rect 17899 19558 17925 19610
rect 17925 19558 17955 19610
rect 17979 19558 17989 19610
rect 17989 19558 18035 19610
rect 18059 19558 18105 19610
rect 18105 19558 18115 19610
rect 18139 19558 18169 19610
rect 18169 19558 18195 19610
rect 17899 19556 17955 19558
rect 17979 19556 18035 19558
rect 18059 19556 18115 19558
rect 18139 19556 18195 19558
rect 17899 18522 17955 18524
rect 17979 18522 18035 18524
rect 18059 18522 18115 18524
rect 18139 18522 18195 18524
rect 17899 18470 17925 18522
rect 17925 18470 17955 18522
rect 17979 18470 17989 18522
rect 17989 18470 18035 18522
rect 18059 18470 18105 18522
rect 18105 18470 18115 18522
rect 18139 18470 18169 18522
rect 18169 18470 18195 18522
rect 17899 18468 17955 18470
rect 17979 18468 18035 18470
rect 18059 18468 18115 18470
rect 18139 18468 18195 18470
rect 17899 17434 17955 17436
rect 17979 17434 18035 17436
rect 18059 17434 18115 17436
rect 18139 17434 18195 17436
rect 17899 17382 17925 17434
rect 17925 17382 17955 17434
rect 17979 17382 17989 17434
rect 17989 17382 18035 17434
rect 18059 17382 18105 17434
rect 18105 17382 18115 17434
rect 18139 17382 18169 17434
rect 18169 17382 18195 17434
rect 17899 17380 17955 17382
rect 17979 17380 18035 17382
rect 18059 17380 18115 17382
rect 18139 17380 18195 17382
rect 17899 16346 17955 16348
rect 17979 16346 18035 16348
rect 18059 16346 18115 16348
rect 18139 16346 18195 16348
rect 17899 16294 17925 16346
rect 17925 16294 17955 16346
rect 17979 16294 17989 16346
rect 17989 16294 18035 16346
rect 18059 16294 18105 16346
rect 18105 16294 18115 16346
rect 18139 16294 18169 16346
rect 18169 16294 18195 16346
rect 17899 16292 17955 16294
rect 17979 16292 18035 16294
rect 18059 16292 18115 16294
rect 18139 16292 18195 16294
rect 17899 15258 17955 15260
rect 17979 15258 18035 15260
rect 18059 15258 18115 15260
rect 18139 15258 18195 15260
rect 17899 15206 17925 15258
rect 17925 15206 17955 15258
rect 17979 15206 17989 15258
rect 17989 15206 18035 15258
rect 18059 15206 18105 15258
rect 18105 15206 18115 15258
rect 18139 15206 18169 15258
rect 18169 15206 18195 15258
rect 17899 15204 17955 15206
rect 17979 15204 18035 15206
rect 18059 15204 18115 15206
rect 18139 15204 18195 15206
rect 19246 14728 19302 14784
rect 17899 14170 17955 14172
rect 17979 14170 18035 14172
rect 18059 14170 18115 14172
rect 18139 14170 18195 14172
rect 17899 14118 17925 14170
rect 17925 14118 17955 14170
rect 17979 14118 17989 14170
rect 17989 14118 18035 14170
rect 18059 14118 18105 14170
rect 18105 14118 18115 14170
rect 18139 14118 18169 14170
rect 18169 14118 18195 14170
rect 17899 14116 17955 14118
rect 17979 14116 18035 14118
rect 18059 14116 18115 14118
rect 18139 14116 18195 14118
rect 17899 13082 17955 13084
rect 17979 13082 18035 13084
rect 18059 13082 18115 13084
rect 18139 13082 18195 13084
rect 17899 13030 17925 13082
rect 17925 13030 17955 13082
rect 17979 13030 17989 13082
rect 17989 13030 18035 13082
rect 18059 13030 18105 13082
rect 18105 13030 18115 13082
rect 18139 13030 18169 13082
rect 18169 13030 18195 13082
rect 17899 13028 17955 13030
rect 17979 13028 18035 13030
rect 18059 13028 18115 13030
rect 18139 13028 18195 13030
rect 17899 11994 17955 11996
rect 17979 11994 18035 11996
rect 18059 11994 18115 11996
rect 18139 11994 18195 11996
rect 17899 11942 17925 11994
rect 17925 11942 17955 11994
rect 17979 11942 17989 11994
rect 17989 11942 18035 11994
rect 18059 11942 18105 11994
rect 18105 11942 18115 11994
rect 18139 11942 18169 11994
rect 18169 11942 18195 11994
rect 17899 11940 17955 11942
rect 17979 11940 18035 11942
rect 18059 11940 18115 11942
rect 18139 11940 18195 11942
rect 17899 10906 17955 10908
rect 17979 10906 18035 10908
rect 18059 10906 18115 10908
rect 18139 10906 18195 10908
rect 17899 10854 17925 10906
rect 17925 10854 17955 10906
rect 17979 10854 17989 10906
rect 17989 10854 18035 10906
rect 18059 10854 18105 10906
rect 18105 10854 18115 10906
rect 18139 10854 18169 10906
rect 18169 10854 18195 10906
rect 17899 10852 17955 10854
rect 17979 10852 18035 10854
rect 18059 10852 18115 10854
rect 18139 10852 18195 10854
rect 17899 9818 17955 9820
rect 17979 9818 18035 9820
rect 18059 9818 18115 9820
rect 18139 9818 18195 9820
rect 17899 9766 17925 9818
rect 17925 9766 17955 9818
rect 17979 9766 17989 9818
rect 17989 9766 18035 9818
rect 18059 9766 18105 9818
rect 18105 9766 18115 9818
rect 18139 9766 18169 9818
rect 18169 9766 18195 9818
rect 17899 9764 17955 9766
rect 17979 9764 18035 9766
rect 18059 9764 18115 9766
rect 18139 9764 18195 9766
rect 17899 8730 17955 8732
rect 17979 8730 18035 8732
rect 18059 8730 18115 8732
rect 18139 8730 18195 8732
rect 17899 8678 17925 8730
rect 17925 8678 17955 8730
rect 17979 8678 17989 8730
rect 17989 8678 18035 8730
rect 18059 8678 18105 8730
rect 18105 8678 18115 8730
rect 18139 8678 18169 8730
rect 18169 8678 18195 8730
rect 17899 8676 17955 8678
rect 17979 8676 18035 8678
rect 18059 8676 18115 8678
rect 18139 8676 18195 8678
rect 17899 7642 17955 7644
rect 17979 7642 18035 7644
rect 18059 7642 18115 7644
rect 18139 7642 18195 7644
rect 17899 7590 17925 7642
rect 17925 7590 17955 7642
rect 17979 7590 17989 7642
rect 17989 7590 18035 7642
rect 18059 7590 18105 7642
rect 18105 7590 18115 7642
rect 18139 7590 18169 7642
rect 18169 7590 18195 7642
rect 17899 7588 17955 7590
rect 17979 7588 18035 7590
rect 18059 7588 18115 7590
rect 18139 7588 18195 7590
rect 17899 6554 17955 6556
rect 17979 6554 18035 6556
rect 18059 6554 18115 6556
rect 18139 6554 18195 6556
rect 17899 6502 17925 6554
rect 17925 6502 17955 6554
rect 17979 6502 17989 6554
rect 17989 6502 18035 6554
rect 18059 6502 18105 6554
rect 18105 6502 18115 6554
rect 18139 6502 18169 6554
rect 18169 6502 18195 6554
rect 17899 6500 17955 6502
rect 17979 6500 18035 6502
rect 18059 6500 18115 6502
rect 18139 6500 18195 6502
rect 18326 5480 18382 5536
rect 17899 5466 17955 5468
rect 17979 5466 18035 5468
rect 18059 5466 18115 5468
rect 18139 5466 18195 5468
rect 17899 5414 17925 5466
rect 17925 5414 17955 5466
rect 17979 5414 17989 5466
rect 17989 5414 18035 5466
rect 18059 5414 18105 5466
rect 18105 5414 18115 5466
rect 18139 5414 18169 5466
rect 18169 5414 18195 5466
rect 17899 5412 17955 5414
rect 17979 5412 18035 5414
rect 18059 5412 18115 5414
rect 18139 5412 18195 5414
rect 17899 4378 17955 4380
rect 17979 4378 18035 4380
rect 18059 4378 18115 4380
rect 18139 4378 18195 4380
rect 17899 4326 17925 4378
rect 17925 4326 17955 4378
rect 17979 4326 17989 4378
rect 17989 4326 18035 4378
rect 18059 4326 18105 4378
rect 18105 4326 18115 4378
rect 18139 4326 18169 4378
rect 18169 4326 18195 4378
rect 17899 4324 17955 4326
rect 17979 4324 18035 4326
rect 18059 4324 18115 4326
rect 18139 4324 18195 4326
rect 17899 3290 17955 3292
rect 17979 3290 18035 3292
rect 18059 3290 18115 3292
rect 18139 3290 18195 3292
rect 17899 3238 17925 3290
rect 17925 3238 17955 3290
rect 17979 3238 17989 3290
rect 17989 3238 18035 3290
rect 18059 3238 18105 3290
rect 18105 3238 18115 3290
rect 18139 3238 18169 3290
rect 18169 3238 18195 3290
rect 17899 3236 17955 3238
rect 17979 3236 18035 3238
rect 18059 3236 18115 3238
rect 18139 3236 18195 3238
rect 17899 2202 17955 2204
rect 17979 2202 18035 2204
rect 18059 2202 18115 2204
rect 18139 2202 18195 2204
rect 17899 2150 17925 2202
rect 17925 2150 17955 2202
rect 17979 2150 17989 2202
rect 17989 2150 18035 2202
rect 18059 2150 18105 2202
rect 18105 2150 18115 2202
rect 18139 2150 18169 2202
rect 18169 2150 18195 2202
rect 17899 2148 17955 2150
rect 17979 2148 18035 2150
rect 18059 2148 18115 2150
rect 18139 2148 18195 2150
<< metal3 >>
rect 7721 22336 8041 22337
rect 7721 22272 7729 22336
rect 7793 22272 7809 22336
rect 7873 22272 7889 22336
rect 7953 22272 7969 22336
rect 8033 22272 8041 22336
rect 7721 22271 8041 22272
rect 14498 22336 14818 22337
rect 14498 22272 14506 22336
rect 14570 22272 14586 22336
rect 14650 22272 14666 22336
rect 14730 22272 14746 22336
rect 14810 22272 14818 22336
rect 14498 22271 14818 22272
rect 4332 21792 4652 21793
rect 4332 21728 4340 21792
rect 4404 21728 4420 21792
rect 4484 21728 4500 21792
rect 4564 21728 4580 21792
rect 4644 21728 4652 21792
rect 4332 21727 4652 21728
rect 11110 21792 11430 21793
rect 11110 21728 11118 21792
rect 11182 21728 11198 21792
rect 11262 21728 11278 21792
rect 11342 21728 11358 21792
rect 11422 21728 11430 21792
rect 11110 21727 11430 21728
rect 17887 21792 18207 21793
rect 17887 21728 17895 21792
rect 17959 21728 17975 21792
rect 18039 21728 18055 21792
rect 18119 21728 18135 21792
rect 18199 21728 18207 21792
rect 17887 21727 18207 21728
rect 7721 21248 8041 21249
rect 7721 21184 7729 21248
rect 7793 21184 7809 21248
rect 7873 21184 7889 21248
rect 7953 21184 7969 21248
rect 8033 21184 8041 21248
rect 7721 21183 8041 21184
rect 14498 21248 14818 21249
rect 14498 21184 14506 21248
rect 14570 21184 14586 21248
rect 14650 21184 14666 21248
rect 14730 21184 14746 21248
rect 14810 21184 14818 21248
rect 14498 21183 14818 21184
rect 4332 20704 4652 20705
rect 4332 20640 4340 20704
rect 4404 20640 4420 20704
rect 4484 20640 4500 20704
rect 4564 20640 4580 20704
rect 4644 20640 4652 20704
rect 4332 20639 4652 20640
rect 11110 20704 11430 20705
rect 11110 20640 11118 20704
rect 11182 20640 11198 20704
rect 11262 20640 11278 20704
rect 11342 20640 11358 20704
rect 11422 20640 11430 20704
rect 11110 20639 11430 20640
rect 17887 20704 18207 20705
rect 17887 20640 17895 20704
rect 17959 20640 17975 20704
rect 18039 20640 18055 20704
rect 18119 20640 18135 20704
rect 18199 20640 18207 20704
rect 17887 20639 18207 20640
rect 7721 20160 8041 20161
rect 7721 20096 7729 20160
rect 7793 20096 7809 20160
rect 7873 20096 7889 20160
rect 7953 20096 7969 20160
rect 8033 20096 8041 20160
rect 7721 20095 8041 20096
rect 14498 20160 14818 20161
rect 14498 20096 14506 20160
rect 14570 20096 14586 20160
rect 14650 20096 14666 20160
rect 14730 20096 14746 20160
rect 14810 20096 14818 20160
rect 14498 20095 14818 20096
rect 4332 19616 4652 19617
rect 4332 19552 4340 19616
rect 4404 19552 4420 19616
rect 4484 19552 4500 19616
rect 4564 19552 4580 19616
rect 4644 19552 4652 19616
rect 4332 19551 4652 19552
rect 11110 19616 11430 19617
rect 11110 19552 11118 19616
rect 11182 19552 11198 19616
rect 11262 19552 11278 19616
rect 11342 19552 11358 19616
rect 11422 19552 11430 19616
rect 11110 19551 11430 19552
rect 17887 19616 18207 19617
rect 17887 19552 17895 19616
rect 17959 19552 17975 19616
rect 18039 19552 18055 19616
rect 18119 19552 18135 19616
rect 18199 19552 18207 19616
rect 17887 19551 18207 19552
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 7721 19072 8041 19073
rect 7721 19008 7729 19072
rect 7793 19008 7809 19072
rect 7873 19008 7889 19072
rect 7953 19008 7969 19072
rect 8033 19008 8041 19072
rect 7721 19007 8041 19008
rect 14498 19072 14818 19073
rect 14498 19008 14506 19072
rect 14570 19008 14586 19072
rect 14650 19008 14666 19072
rect 14730 19008 14746 19072
rect 14810 19008 14818 19072
rect 14498 19007 14818 19008
rect 4332 18528 4652 18529
rect 4332 18464 4340 18528
rect 4404 18464 4420 18528
rect 4484 18464 4500 18528
rect 4564 18464 4580 18528
rect 4644 18464 4652 18528
rect 4332 18463 4652 18464
rect 11110 18528 11430 18529
rect 11110 18464 11118 18528
rect 11182 18464 11198 18528
rect 11262 18464 11278 18528
rect 11342 18464 11358 18528
rect 11422 18464 11430 18528
rect 11110 18463 11430 18464
rect 17887 18528 18207 18529
rect 17887 18464 17895 18528
rect 17959 18464 17975 18528
rect 18039 18464 18055 18528
rect 18119 18464 18135 18528
rect 18199 18464 18207 18528
rect 17887 18463 18207 18464
rect 7721 17984 8041 17985
rect 7721 17920 7729 17984
rect 7793 17920 7809 17984
rect 7873 17920 7889 17984
rect 7953 17920 7969 17984
rect 8033 17920 8041 17984
rect 7721 17919 8041 17920
rect 14498 17984 14818 17985
rect 14498 17920 14506 17984
rect 14570 17920 14586 17984
rect 14650 17920 14666 17984
rect 14730 17920 14746 17984
rect 14810 17920 14818 17984
rect 14498 17919 14818 17920
rect 4332 17440 4652 17441
rect 4332 17376 4340 17440
rect 4404 17376 4420 17440
rect 4484 17376 4500 17440
rect 4564 17376 4580 17440
rect 4644 17376 4652 17440
rect 4332 17375 4652 17376
rect 11110 17440 11430 17441
rect 11110 17376 11118 17440
rect 11182 17376 11198 17440
rect 11262 17376 11278 17440
rect 11342 17376 11358 17440
rect 11422 17376 11430 17440
rect 11110 17375 11430 17376
rect 17887 17440 18207 17441
rect 17887 17376 17895 17440
rect 17959 17376 17975 17440
rect 18039 17376 18055 17440
rect 18119 17376 18135 17440
rect 18199 17376 18207 17440
rect 17887 17375 18207 17376
rect 7721 16896 8041 16897
rect 7721 16832 7729 16896
rect 7793 16832 7809 16896
rect 7873 16832 7889 16896
rect 7953 16832 7969 16896
rect 8033 16832 8041 16896
rect 7721 16831 8041 16832
rect 14498 16896 14818 16897
rect 14498 16832 14506 16896
rect 14570 16832 14586 16896
rect 14650 16832 14666 16896
rect 14730 16832 14746 16896
rect 14810 16832 14818 16896
rect 14498 16831 14818 16832
rect 4332 16352 4652 16353
rect 4332 16288 4340 16352
rect 4404 16288 4420 16352
rect 4484 16288 4500 16352
rect 4564 16288 4580 16352
rect 4644 16288 4652 16352
rect 4332 16287 4652 16288
rect 11110 16352 11430 16353
rect 11110 16288 11118 16352
rect 11182 16288 11198 16352
rect 11262 16288 11278 16352
rect 11342 16288 11358 16352
rect 11422 16288 11430 16352
rect 11110 16287 11430 16288
rect 17887 16352 18207 16353
rect 17887 16288 17895 16352
rect 17959 16288 17975 16352
rect 18039 16288 18055 16352
rect 18119 16288 18135 16352
rect 18199 16288 18207 16352
rect 17887 16287 18207 16288
rect 7721 15808 8041 15809
rect 7721 15744 7729 15808
rect 7793 15744 7809 15808
rect 7873 15744 7889 15808
rect 7953 15744 7969 15808
rect 8033 15744 8041 15808
rect 7721 15743 8041 15744
rect 14498 15808 14818 15809
rect 14498 15744 14506 15808
rect 14570 15744 14586 15808
rect 14650 15744 14666 15808
rect 14730 15744 14746 15808
rect 14810 15744 14818 15808
rect 14498 15743 14818 15744
rect 4332 15264 4652 15265
rect 4332 15200 4340 15264
rect 4404 15200 4420 15264
rect 4484 15200 4500 15264
rect 4564 15200 4580 15264
rect 4644 15200 4652 15264
rect 4332 15199 4652 15200
rect 11110 15264 11430 15265
rect 11110 15200 11118 15264
rect 11182 15200 11198 15264
rect 11262 15200 11278 15264
rect 11342 15200 11358 15264
rect 11422 15200 11430 15264
rect 11110 15199 11430 15200
rect 17887 15264 18207 15265
rect 17887 15200 17895 15264
rect 17959 15200 17975 15264
rect 18039 15200 18055 15264
rect 18119 15200 18135 15264
rect 18199 15200 18207 15264
rect 17887 15199 18207 15200
rect 19241 14786 19307 14789
rect 21789 14786 22589 14816
rect 19241 14784 22589 14786
rect 19241 14728 19246 14784
rect 19302 14728 22589 14784
rect 19241 14726 22589 14728
rect 19241 14723 19307 14726
rect 7721 14720 8041 14721
rect 7721 14656 7729 14720
rect 7793 14656 7809 14720
rect 7873 14656 7889 14720
rect 7953 14656 7969 14720
rect 8033 14656 8041 14720
rect 7721 14655 8041 14656
rect 14498 14720 14818 14721
rect 14498 14656 14506 14720
rect 14570 14656 14586 14720
rect 14650 14656 14666 14720
rect 14730 14656 14746 14720
rect 14810 14656 14818 14720
rect 21789 14696 22589 14726
rect 14498 14655 14818 14656
rect 4332 14176 4652 14177
rect 4332 14112 4340 14176
rect 4404 14112 4420 14176
rect 4484 14112 4500 14176
rect 4564 14112 4580 14176
rect 4644 14112 4652 14176
rect 4332 14111 4652 14112
rect 11110 14176 11430 14177
rect 11110 14112 11118 14176
rect 11182 14112 11198 14176
rect 11262 14112 11278 14176
rect 11342 14112 11358 14176
rect 11422 14112 11430 14176
rect 11110 14111 11430 14112
rect 17887 14176 18207 14177
rect 17887 14112 17895 14176
rect 17959 14112 17975 14176
rect 18039 14112 18055 14176
rect 18119 14112 18135 14176
rect 18199 14112 18207 14176
rect 17887 14111 18207 14112
rect 7721 13632 8041 13633
rect 7721 13568 7729 13632
rect 7793 13568 7809 13632
rect 7873 13568 7889 13632
rect 7953 13568 7969 13632
rect 8033 13568 8041 13632
rect 7721 13567 8041 13568
rect 14498 13632 14818 13633
rect 14498 13568 14506 13632
rect 14570 13568 14586 13632
rect 14650 13568 14666 13632
rect 14730 13568 14746 13632
rect 14810 13568 14818 13632
rect 14498 13567 14818 13568
rect 4332 13088 4652 13089
rect 4332 13024 4340 13088
rect 4404 13024 4420 13088
rect 4484 13024 4500 13088
rect 4564 13024 4580 13088
rect 4644 13024 4652 13088
rect 4332 13023 4652 13024
rect 11110 13088 11430 13089
rect 11110 13024 11118 13088
rect 11182 13024 11198 13088
rect 11262 13024 11278 13088
rect 11342 13024 11358 13088
rect 11422 13024 11430 13088
rect 11110 13023 11430 13024
rect 17887 13088 18207 13089
rect 17887 13024 17895 13088
rect 17959 13024 17975 13088
rect 18039 13024 18055 13088
rect 18119 13024 18135 13088
rect 18199 13024 18207 13088
rect 17887 13023 18207 13024
rect 7721 12544 8041 12545
rect 7721 12480 7729 12544
rect 7793 12480 7809 12544
rect 7873 12480 7889 12544
rect 7953 12480 7969 12544
rect 8033 12480 8041 12544
rect 7721 12479 8041 12480
rect 14498 12544 14818 12545
rect 14498 12480 14506 12544
rect 14570 12480 14586 12544
rect 14650 12480 14666 12544
rect 14730 12480 14746 12544
rect 14810 12480 14818 12544
rect 14498 12479 14818 12480
rect 4332 12000 4652 12001
rect 4332 11936 4340 12000
rect 4404 11936 4420 12000
rect 4484 11936 4500 12000
rect 4564 11936 4580 12000
rect 4644 11936 4652 12000
rect 4332 11935 4652 11936
rect 11110 12000 11430 12001
rect 11110 11936 11118 12000
rect 11182 11936 11198 12000
rect 11262 11936 11278 12000
rect 11342 11936 11358 12000
rect 11422 11936 11430 12000
rect 11110 11935 11430 11936
rect 17887 12000 18207 12001
rect 17887 11936 17895 12000
rect 17959 11936 17975 12000
rect 18039 11936 18055 12000
rect 18119 11936 18135 12000
rect 18199 11936 18207 12000
rect 17887 11935 18207 11936
rect 7721 11456 8041 11457
rect 7721 11392 7729 11456
rect 7793 11392 7809 11456
rect 7873 11392 7889 11456
rect 7953 11392 7969 11456
rect 8033 11392 8041 11456
rect 7721 11391 8041 11392
rect 14498 11456 14818 11457
rect 14498 11392 14506 11456
rect 14570 11392 14586 11456
rect 14650 11392 14666 11456
rect 14730 11392 14746 11456
rect 14810 11392 14818 11456
rect 14498 11391 14818 11392
rect 4332 10912 4652 10913
rect 4332 10848 4340 10912
rect 4404 10848 4420 10912
rect 4484 10848 4500 10912
rect 4564 10848 4580 10912
rect 4644 10848 4652 10912
rect 4332 10847 4652 10848
rect 11110 10912 11430 10913
rect 11110 10848 11118 10912
rect 11182 10848 11198 10912
rect 11262 10848 11278 10912
rect 11342 10848 11358 10912
rect 11422 10848 11430 10912
rect 11110 10847 11430 10848
rect 17887 10912 18207 10913
rect 17887 10848 17895 10912
rect 17959 10848 17975 10912
rect 18039 10848 18055 10912
rect 18119 10848 18135 10912
rect 18199 10848 18207 10912
rect 17887 10847 18207 10848
rect 7721 10368 8041 10369
rect 7721 10304 7729 10368
rect 7793 10304 7809 10368
rect 7873 10304 7889 10368
rect 7953 10304 7969 10368
rect 8033 10304 8041 10368
rect 7721 10303 8041 10304
rect 14498 10368 14818 10369
rect 14498 10304 14506 10368
rect 14570 10304 14586 10368
rect 14650 10304 14666 10368
rect 14730 10304 14746 10368
rect 14810 10304 14818 10368
rect 14498 10303 14818 10304
rect 0 9890 800 9920
rect 4061 9890 4127 9893
rect 0 9888 4127 9890
rect 0 9832 4066 9888
rect 4122 9832 4127 9888
rect 0 9830 4127 9832
rect 0 9800 800 9830
rect 4061 9827 4127 9830
rect 4332 9824 4652 9825
rect 4332 9760 4340 9824
rect 4404 9760 4420 9824
rect 4484 9760 4500 9824
rect 4564 9760 4580 9824
rect 4644 9760 4652 9824
rect 4332 9759 4652 9760
rect 11110 9824 11430 9825
rect 11110 9760 11118 9824
rect 11182 9760 11198 9824
rect 11262 9760 11278 9824
rect 11342 9760 11358 9824
rect 11422 9760 11430 9824
rect 11110 9759 11430 9760
rect 17887 9824 18207 9825
rect 17887 9760 17895 9824
rect 17959 9760 17975 9824
rect 18039 9760 18055 9824
rect 18119 9760 18135 9824
rect 18199 9760 18207 9824
rect 17887 9759 18207 9760
rect 4797 9754 4863 9757
rect 5349 9754 5415 9757
rect 4797 9752 5415 9754
rect 4797 9696 4802 9752
rect 4858 9696 5354 9752
rect 5410 9696 5415 9752
rect 4797 9694 5415 9696
rect 4797 9691 4863 9694
rect 5349 9691 5415 9694
rect 13261 9754 13327 9757
rect 13261 9752 15394 9754
rect 13261 9696 13266 9752
rect 13322 9696 15394 9752
rect 13261 9694 15394 9696
rect 13261 9691 13327 9694
rect 12617 9652 12683 9655
rect 12617 9650 12818 9652
rect 12617 9594 12622 9650
rect 12678 9618 12818 9650
rect 12985 9618 13051 9621
rect 12678 9616 13051 9618
rect 12678 9594 12990 9616
rect 12617 9592 12990 9594
rect 12617 9589 12683 9592
rect 12758 9560 12990 9592
rect 13046 9560 13051 9616
rect 12758 9558 13051 9560
rect 15334 9618 15394 9694
rect 15837 9618 15903 9621
rect 15334 9616 15903 9618
rect 15334 9560 15842 9616
rect 15898 9560 15903 9616
rect 15334 9558 15903 9560
rect 12985 9555 13051 9558
rect 15837 9555 15903 9558
rect 7721 9280 8041 9281
rect 7721 9216 7729 9280
rect 7793 9216 7809 9280
rect 7873 9216 7889 9280
rect 7953 9216 7969 9280
rect 8033 9216 8041 9280
rect 7721 9215 8041 9216
rect 14498 9280 14818 9281
rect 14498 9216 14506 9280
rect 14570 9216 14586 9280
rect 14650 9216 14666 9280
rect 14730 9216 14746 9280
rect 14810 9216 14818 9280
rect 14498 9215 14818 9216
rect 4332 8736 4652 8737
rect 4332 8672 4340 8736
rect 4404 8672 4420 8736
rect 4484 8672 4500 8736
rect 4564 8672 4580 8736
rect 4644 8672 4652 8736
rect 4332 8671 4652 8672
rect 11110 8736 11430 8737
rect 11110 8672 11118 8736
rect 11182 8672 11198 8736
rect 11262 8672 11278 8736
rect 11342 8672 11358 8736
rect 11422 8672 11430 8736
rect 11110 8671 11430 8672
rect 17887 8736 18207 8737
rect 17887 8672 17895 8736
rect 17959 8672 17975 8736
rect 18039 8672 18055 8736
rect 18119 8672 18135 8736
rect 18199 8672 18207 8736
rect 17887 8671 18207 8672
rect 12893 8530 12959 8533
rect 15745 8530 15811 8533
rect 12893 8528 15811 8530
rect 12893 8472 12898 8528
rect 12954 8472 15750 8528
rect 15806 8472 15811 8528
rect 12893 8470 15811 8472
rect 12893 8467 12959 8470
rect 15745 8467 15811 8470
rect 7721 8192 8041 8193
rect 7721 8128 7729 8192
rect 7793 8128 7809 8192
rect 7873 8128 7889 8192
rect 7953 8128 7969 8192
rect 8033 8128 8041 8192
rect 7721 8127 8041 8128
rect 14498 8192 14818 8193
rect 14498 8128 14506 8192
rect 14570 8128 14586 8192
rect 14650 8128 14666 8192
rect 14730 8128 14746 8192
rect 14810 8128 14818 8192
rect 14498 8127 14818 8128
rect 4332 7648 4652 7649
rect 4332 7584 4340 7648
rect 4404 7584 4420 7648
rect 4484 7584 4500 7648
rect 4564 7584 4580 7648
rect 4644 7584 4652 7648
rect 4332 7583 4652 7584
rect 11110 7648 11430 7649
rect 11110 7584 11118 7648
rect 11182 7584 11198 7648
rect 11262 7584 11278 7648
rect 11342 7584 11358 7648
rect 11422 7584 11430 7648
rect 11110 7583 11430 7584
rect 17887 7648 18207 7649
rect 17887 7584 17895 7648
rect 17959 7584 17975 7648
rect 18039 7584 18055 7648
rect 18119 7584 18135 7648
rect 18199 7584 18207 7648
rect 17887 7583 18207 7584
rect 7721 7104 8041 7105
rect 7721 7040 7729 7104
rect 7793 7040 7809 7104
rect 7873 7040 7889 7104
rect 7953 7040 7969 7104
rect 8033 7040 8041 7104
rect 7721 7039 8041 7040
rect 14498 7104 14818 7105
rect 14498 7040 14506 7104
rect 14570 7040 14586 7104
rect 14650 7040 14666 7104
rect 14730 7040 14746 7104
rect 14810 7040 14818 7104
rect 14498 7039 14818 7040
rect 4332 6560 4652 6561
rect 4332 6496 4340 6560
rect 4404 6496 4420 6560
rect 4484 6496 4500 6560
rect 4564 6496 4580 6560
rect 4644 6496 4652 6560
rect 4332 6495 4652 6496
rect 11110 6560 11430 6561
rect 11110 6496 11118 6560
rect 11182 6496 11198 6560
rect 11262 6496 11278 6560
rect 11342 6496 11358 6560
rect 11422 6496 11430 6560
rect 11110 6495 11430 6496
rect 17887 6560 18207 6561
rect 17887 6496 17895 6560
rect 17959 6496 17975 6560
rect 18039 6496 18055 6560
rect 18119 6496 18135 6560
rect 18199 6496 18207 6560
rect 17887 6495 18207 6496
rect 7721 6016 8041 6017
rect 7721 5952 7729 6016
rect 7793 5952 7809 6016
rect 7873 5952 7889 6016
rect 7953 5952 7969 6016
rect 8033 5952 8041 6016
rect 7721 5951 8041 5952
rect 14498 6016 14818 6017
rect 14498 5952 14506 6016
rect 14570 5952 14586 6016
rect 14650 5952 14666 6016
rect 14730 5952 14746 6016
rect 14810 5952 14818 6016
rect 14498 5951 14818 5952
rect 18321 5538 18387 5541
rect 21789 5538 22589 5568
rect 18321 5536 22589 5538
rect 18321 5480 18326 5536
rect 18382 5480 22589 5536
rect 18321 5478 22589 5480
rect 18321 5475 18387 5478
rect 4332 5472 4652 5473
rect 4332 5408 4340 5472
rect 4404 5408 4420 5472
rect 4484 5408 4500 5472
rect 4564 5408 4580 5472
rect 4644 5408 4652 5472
rect 4332 5407 4652 5408
rect 11110 5472 11430 5473
rect 11110 5408 11118 5472
rect 11182 5408 11198 5472
rect 11262 5408 11278 5472
rect 11342 5408 11358 5472
rect 11422 5408 11430 5472
rect 11110 5407 11430 5408
rect 17887 5472 18207 5473
rect 17887 5408 17895 5472
rect 17959 5408 17975 5472
rect 18039 5408 18055 5472
rect 18119 5408 18135 5472
rect 18199 5408 18207 5472
rect 21789 5448 22589 5478
rect 17887 5407 18207 5408
rect 7721 4928 8041 4929
rect 7721 4864 7729 4928
rect 7793 4864 7809 4928
rect 7873 4864 7889 4928
rect 7953 4864 7969 4928
rect 8033 4864 8041 4928
rect 7721 4863 8041 4864
rect 14498 4928 14818 4929
rect 14498 4864 14506 4928
rect 14570 4864 14586 4928
rect 14650 4864 14666 4928
rect 14730 4864 14746 4928
rect 14810 4864 14818 4928
rect 14498 4863 14818 4864
rect 4332 4384 4652 4385
rect 4332 4320 4340 4384
rect 4404 4320 4420 4384
rect 4484 4320 4500 4384
rect 4564 4320 4580 4384
rect 4644 4320 4652 4384
rect 4332 4319 4652 4320
rect 11110 4384 11430 4385
rect 11110 4320 11118 4384
rect 11182 4320 11198 4384
rect 11262 4320 11278 4384
rect 11342 4320 11358 4384
rect 11422 4320 11430 4384
rect 11110 4319 11430 4320
rect 17887 4384 18207 4385
rect 17887 4320 17895 4384
rect 17959 4320 17975 4384
rect 18039 4320 18055 4384
rect 18119 4320 18135 4384
rect 18199 4320 18207 4384
rect 17887 4319 18207 4320
rect 7721 3840 8041 3841
rect 7721 3776 7729 3840
rect 7793 3776 7809 3840
rect 7873 3776 7889 3840
rect 7953 3776 7969 3840
rect 8033 3776 8041 3840
rect 7721 3775 8041 3776
rect 14498 3840 14818 3841
rect 14498 3776 14506 3840
rect 14570 3776 14586 3840
rect 14650 3776 14666 3840
rect 14730 3776 14746 3840
rect 14810 3776 14818 3840
rect 14498 3775 14818 3776
rect 4332 3296 4652 3297
rect 4332 3232 4340 3296
rect 4404 3232 4420 3296
rect 4484 3232 4500 3296
rect 4564 3232 4580 3296
rect 4644 3232 4652 3296
rect 4332 3231 4652 3232
rect 11110 3296 11430 3297
rect 11110 3232 11118 3296
rect 11182 3232 11198 3296
rect 11262 3232 11278 3296
rect 11342 3232 11358 3296
rect 11422 3232 11430 3296
rect 11110 3231 11430 3232
rect 17887 3296 18207 3297
rect 17887 3232 17895 3296
rect 17959 3232 17975 3296
rect 18039 3232 18055 3296
rect 18119 3232 18135 3296
rect 18199 3232 18207 3296
rect 17887 3231 18207 3232
rect 7721 2752 8041 2753
rect 7721 2688 7729 2752
rect 7793 2688 7809 2752
rect 7873 2688 7889 2752
rect 7953 2688 7969 2752
rect 8033 2688 8041 2752
rect 7721 2687 8041 2688
rect 14498 2752 14818 2753
rect 14498 2688 14506 2752
rect 14570 2688 14586 2752
rect 14650 2688 14666 2752
rect 14730 2688 14746 2752
rect 14810 2688 14818 2752
rect 14498 2687 14818 2688
rect 4332 2208 4652 2209
rect 4332 2144 4340 2208
rect 4404 2144 4420 2208
rect 4484 2144 4500 2208
rect 4564 2144 4580 2208
rect 4644 2144 4652 2208
rect 4332 2143 4652 2144
rect 11110 2208 11430 2209
rect 11110 2144 11118 2208
rect 11182 2144 11198 2208
rect 11262 2144 11278 2208
rect 11342 2144 11358 2208
rect 11422 2144 11430 2208
rect 11110 2143 11430 2144
rect 17887 2208 18207 2209
rect 17887 2144 17895 2208
rect 17959 2144 17975 2208
rect 18039 2144 18055 2208
rect 18119 2144 18135 2208
rect 18199 2144 18207 2208
rect 17887 2143 18207 2144
<< via3 >>
rect 7729 22332 7793 22336
rect 7729 22276 7733 22332
rect 7733 22276 7789 22332
rect 7789 22276 7793 22332
rect 7729 22272 7793 22276
rect 7809 22332 7873 22336
rect 7809 22276 7813 22332
rect 7813 22276 7869 22332
rect 7869 22276 7873 22332
rect 7809 22272 7873 22276
rect 7889 22332 7953 22336
rect 7889 22276 7893 22332
rect 7893 22276 7949 22332
rect 7949 22276 7953 22332
rect 7889 22272 7953 22276
rect 7969 22332 8033 22336
rect 7969 22276 7973 22332
rect 7973 22276 8029 22332
rect 8029 22276 8033 22332
rect 7969 22272 8033 22276
rect 14506 22332 14570 22336
rect 14506 22276 14510 22332
rect 14510 22276 14566 22332
rect 14566 22276 14570 22332
rect 14506 22272 14570 22276
rect 14586 22332 14650 22336
rect 14586 22276 14590 22332
rect 14590 22276 14646 22332
rect 14646 22276 14650 22332
rect 14586 22272 14650 22276
rect 14666 22332 14730 22336
rect 14666 22276 14670 22332
rect 14670 22276 14726 22332
rect 14726 22276 14730 22332
rect 14666 22272 14730 22276
rect 14746 22332 14810 22336
rect 14746 22276 14750 22332
rect 14750 22276 14806 22332
rect 14806 22276 14810 22332
rect 14746 22272 14810 22276
rect 4340 21788 4404 21792
rect 4340 21732 4344 21788
rect 4344 21732 4400 21788
rect 4400 21732 4404 21788
rect 4340 21728 4404 21732
rect 4420 21788 4484 21792
rect 4420 21732 4424 21788
rect 4424 21732 4480 21788
rect 4480 21732 4484 21788
rect 4420 21728 4484 21732
rect 4500 21788 4564 21792
rect 4500 21732 4504 21788
rect 4504 21732 4560 21788
rect 4560 21732 4564 21788
rect 4500 21728 4564 21732
rect 4580 21788 4644 21792
rect 4580 21732 4584 21788
rect 4584 21732 4640 21788
rect 4640 21732 4644 21788
rect 4580 21728 4644 21732
rect 11118 21788 11182 21792
rect 11118 21732 11122 21788
rect 11122 21732 11178 21788
rect 11178 21732 11182 21788
rect 11118 21728 11182 21732
rect 11198 21788 11262 21792
rect 11198 21732 11202 21788
rect 11202 21732 11258 21788
rect 11258 21732 11262 21788
rect 11198 21728 11262 21732
rect 11278 21788 11342 21792
rect 11278 21732 11282 21788
rect 11282 21732 11338 21788
rect 11338 21732 11342 21788
rect 11278 21728 11342 21732
rect 11358 21788 11422 21792
rect 11358 21732 11362 21788
rect 11362 21732 11418 21788
rect 11418 21732 11422 21788
rect 11358 21728 11422 21732
rect 17895 21788 17959 21792
rect 17895 21732 17899 21788
rect 17899 21732 17955 21788
rect 17955 21732 17959 21788
rect 17895 21728 17959 21732
rect 17975 21788 18039 21792
rect 17975 21732 17979 21788
rect 17979 21732 18035 21788
rect 18035 21732 18039 21788
rect 17975 21728 18039 21732
rect 18055 21788 18119 21792
rect 18055 21732 18059 21788
rect 18059 21732 18115 21788
rect 18115 21732 18119 21788
rect 18055 21728 18119 21732
rect 18135 21788 18199 21792
rect 18135 21732 18139 21788
rect 18139 21732 18195 21788
rect 18195 21732 18199 21788
rect 18135 21728 18199 21732
rect 7729 21244 7793 21248
rect 7729 21188 7733 21244
rect 7733 21188 7789 21244
rect 7789 21188 7793 21244
rect 7729 21184 7793 21188
rect 7809 21244 7873 21248
rect 7809 21188 7813 21244
rect 7813 21188 7869 21244
rect 7869 21188 7873 21244
rect 7809 21184 7873 21188
rect 7889 21244 7953 21248
rect 7889 21188 7893 21244
rect 7893 21188 7949 21244
rect 7949 21188 7953 21244
rect 7889 21184 7953 21188
rect 7969 21244 8033 21248
rect 7969 21188 7973 21244
rect 7973 21188 8029 21244
rect 8029 21188 8033 21244
rect 7969 21184 8033 21188
rect 14506 21244 14570 21248
rect 14506 21188 14510 21244
rect 14510 21188 14566 21244
rect 14566 21188 14570 21244
rect 14506 21184 14570 21188
rect 14586 21244 14650 21248
rect 14586 21188 14590 21244
rect 14590 21188 14646 21244
rect 14646 21188 14650 21244
rect 14586 21184 14650 21188
rect 14666 21244 14730 21248
rect 14666 21188 14670 21244
rect 14670 21188 14726 21244
rect 14726 21188 14730 21244
rect 14666 21184 14730 21188
rect 14746 21244 14810 21248
rect 14746 21188 14750 21244
rect 14750 21188 14806 21244
rect 14806 21188 14810 21244
rect 14746 21184 14810 21188
rect 4340 20700 4404 20704
rect 4340 20644 4344 20700
rect 4344 20644 4400 20700
rect 4400 20644 4404 20700
rect 4340 20640 4404 20644
rect 4420 20700 4484 20704
rect 4420 20644 4424 20700
rect 4424 20644 4480 20700
rect 4480 20644 4484 20700
rect 4420 20640 4484 20644
rect 4500 20700 4564 20704
rect 4500 20644 4504 20700
rect 4504 20644 4560 20700
rect 4560 20644 4564 20700
rect 4500 20640 4564 20644
rect 4580 20700 4644 20704
rect 4580 20644 4584 20700
rect 4584 20644 4640 20700
rect 4640 20644 4644 20700
rect 4580 20640 4644 20644
rect 11118 20700 11182 20704
rect 11118 20644 11122 20700
rect 11122 20644 11178 20700
rect 11178 20644 11182 20700
rect 11118 20640 11182 20644
rect 11198 20700 11262 20704
rect 11198 20644 11202 20700
rect 11202 20644 11258 20700
rect 11258 20644 11262 20700
rect 11198 20640 11262 20644
rect 11278 20700 11342 20704
rect 11278 20644 11282 20700
rect 11282 20644 11338 20700
rect 11338 20644 11342 20700
rect 11278 20640 11342 20644
rect 11358 20700 11422 20704
rect 11358 20644 11362 20700
rect 11362 20644 11418 20700
rect 11418 20644 11422 20700
rect 11358 20640 11422 20644
rect 17895 20700 17959 20704
rect 17895 20644 17899 20700
rect 17899 20644 17955 20700
rect 17955 20644 17959 20700
rect 17895 20640 17959 20644
rect 17975 20700 18039 20704
rect 17975 20644 17979 20700
rect 17979 20644 18035 20700
rect 18035 20644 18039 20700
rect 17975 20640 18039 20644
rect 18055 20700 18119 20704
rect 18055 20644 18059 20700
rect 18059 20644 18115 20700
rect 18115 20644 18119 20700
rect 18055 20640 18119 20644
rect 18135 20700 18199 20704
rect 18135 20644 18139 20700
rect 18139 20644 18195 20700
rect 18195 20644 18199 20700
rect 18135 20640 18199 20644
rect 7729 20156 7793 20160
rect 7729 20100 7733 20156
rect 7733 20100 7789 20156
rect 7789 20100 7793 20156
rect 7729 20096 7793 20100
rect 7809 20156 7873 20160
rect 7809 20100 7813 20156
rect 7813 20100 7869 20156
rect 7869 20100 7873 20156
rect 7809 20096 7873 20100
rect 7889 20156 7953 20160
rect 7889 20100 7893 20156
rect 7893 20100 7949 20156
rect 7949 20100 7953 20156
rect 7889 20096 7953 20100
rect 7969 20156 8033 20160
rect 7969 20100 7973 20156
rect 7973 20100 8029 20156
rect 8029 20100 8033 20156
rect 7969 20096 8033 20100
rect 14506 20156 14570 20160
rect 14506 20100 14510 20156
rect 14510 20100 14566 20156
rect 14566 20100 14570 20156
rect 14506 20096 14570 20100
rect 14586 20156 14650 20160
rect 14586 20100 14590 20156
rect 14590 20100 14646 20156
rect 14646 20100 14650 20156
rect 14586 20096 14650 20100
rect 14666 20156 14730 20160
rect 14666 20100 14670 20156
rect 14670 20100 14726 20156
rect 14726 20100 14730 20156
rect 14666 20096 14730 20100
rect 14746 20156 14810 20160
rect 14746 20100 14750 20156
rect 14750 20100 14806 20156
rect 14806 20100 14810 20156
rect 14746 20096 14810 20100
rect 4340 19612 4404 19616
rect 4340 19556 4344 19612
rect 4344 19556 4400 19612
rect 4400 19556 4404 19612
rect 4340 19552 4404 19556
rect 4420 19612 4484 19616
rect 4420 19556 4424 19612
rect 4424 19556 4480 19612
rect 4480 19556 4484 19612
rect 4420 19552 4484 19556
rect 4500 19612 4564 19616
rect 4500 19556 4504 19612
rect 4504 19556 4560 19612
rect 4560 19556 4564 19612
rect 4500 19552 4564 19556
rect 4580 19612 4644 19616
rect 4580 19556 4584 19612
rect 4584 19556 4640 19612
rect 4640 19556 4644 19612
rect 4580 19552 4644 19556
rect 11118 19612 11182 19616
rect 11118 19556 11122 19612
rect 11122 19556 11178 19612
rect 11178 19556 11182 19612
rect 11118 19552 11182 19556
rect 11198 19612 11262 19616
rect 11198 19556 11202 19612
rect 11202 19556 11258 19612
rect 11258 19556 11262 19612
rect 11198 19552 11262 19556
rect 11278 19612 11342 19616
rect 11278 19556 11282 19612
rect 11282 19556 11338 19612
rect 11338 19556 11342 19612
rect 11278 19552 11342 19556
rect 11358 19612 11422 19616
rect 11358 19556 11362 19612
rect 11362 19556 11418 19612
rect 11418 19556 11422 19612
rect 11358 19552 11422 19556
rect 17895 19612 17959 19616
rect 17895 19556 17899 19612
rect 17899 19556 17955 19612
rect 17955 19556 17959 19612
rect 17895 19552 17959 19556
rect 17975 19612 18039 19616
rect 17975 19556 17979 19612
rect 17979 19556 18035 19612
rect 18035 19556 18039 19612
rect 17975 19552 18039 19556
rect 18055 19612 18119 19616
rect 18055 19556 18059 19612
rect 18059 19556 18115 19612
rect 18115 19556 18119 19612
rect 18055 19552 18119 19556
rect 18135 19612 18199 19616
rect 18135 19556 18139 19612
rect 18139 19556 18195 19612
rect 18195 19556 18199 19612
rect 18135 19552 18199 19556
rect 7729 19068 7793 19072
rect 7729 19012 7733 19068
rect 7733 19012 7789 19068
rect 7789 19012 7793 19068
rect 7729 19008 7793 19012
rect 7809 19068 7873 19072
rect 7809 19012 7813 19068
rect 7813 19012 7869 19068
rect 7869 19012 7873 19068
rect 7809 19008 7873 19012
rect 7889 19068 7953 19072
rect 7889 19012 7893 19068
rect 7893 19012 7949 19068
rect 7949 19012 7953 19068
rect 7889 19008 7953 19012
rect 7969 19068 8033 19072
rect 7969 19012 7973 19068
rect 7973 19012 8029 19068
rect 8029 19012 8033 19068
rect 7969 19008 8033 19012
rect 14506 19068 14570 19072
rect 14506 19012 14510 19068
rect 14510 19012 14566 19068
rect 14566 19012 14570 19068
rect 14506 19008 14570 19012
rect 14586 19068 14650 19072
rect 14586 19012 14590 19068
rect 14590 19012 14646 19068
rect 14646 19012 14650 19068
rect 14586 19008 14650 19012
rect 14666 19068 14730 19072
rect 14666 19012 14670 19068
rect 14670 19012 14726 19068
rect 14726 19012 14730 19068
rect 14666 19008 14730 19012
rect 14746 19068 14810 19072
rect 14746 19012 14750 19068
rect 14750 19012 14806 19068
rect 14806 19012 14810 19068
rect 14746 19008 14810 19012
rect 4340 18524 4404 18528
rect 4340 18468 4344 18524
rect 4344 18468 4400 18524
rect 4400 18468 4404 18524
rect 4340 18464 4404 18468
rect 4420 18524 4484 18528
rect 4420 18468 4424 18524
rect 4424 18468 4480 18524
rect 4480 18468 4484 18524
rect 4420 18464 4484 18468
rect 4500 18524 4564 18528
rect 4500 18468 4504 18524
rect 4504 18468 4560 18524
rect 4560 18468 4564 18524
rect 4500 18464 4564 18468
rect 4580 18524 4644 18528
rect 4580 18468 4584 18524
rect 4584 18468 4640 18524
rect 4640 18468 4644 18524
rect 4580 18464 4644 18468
rect 11118 18524 11182 18528
rect 11118 18468 11122 18524
rect 11122 18468 11178 18524
rect 11178 18468 11182 18524
rect 11118 18464 11182 18468
rect 11198 18524 11262 18528
rect 11198 18468 11202 18524
rect 11202 18468 11258 18524
rect 11258 18468 11262 18524
rect 11198 18464 11262 18468
rect 11278 18524 11342 18528
rect 11278 18468 11282 18524
rect 11282 18468 11338 18524
rect 11338 18468 11342 18524
rect 11278 18464 11342 18468
rect 11358 18524 11422 18528
rect 11358 18468 11362 18524
rect 11362 18468 11418 18524
rect 11418 18468 11422 18524
rect 11358 18464 11422 18468
rect 17895 18524 17959 18528
rect 17895 18468 17899 18524
rect 17899 18468 17955 18524
rect 17955 18468 17959 18524
rect 17895 18464 17959 18468
rect 17975 18524 18039 18528
rect 17975 18468 17979 18524
rect 17979 18468 18035 18524
rect 18035 18468 18039 18524
rect 17975 18464 18039 18468
rect 18055 18524 18119 18528
rect 18055 18468 18059 18524
rect 18059 18468 18115 18524
rect 18115 18468 18119 18524
rect 18055 18464 18119 18468
rect 18135 18524 18199 18528
rect 18135 18468 18139 18524
rect 18139 18468 18195 18524
rect 18195 18468 18199 18524
rect 18135 18464 18199 18468
rect 7729 17980 7793 17984
rect 7729 17924 7733 17980
rect 7733 17924 7789 17980
rect 7789 17924 7793 17980
rect 7729 17920 7793 17924
rect 7809 17980 7873 17984
rect 7809 17924 7813 17980
rect 7813 17924 7869 17980
rect 7869 17924 7873 17980
rect 7809 17920 7873 17924
rect 7889 17980 7953 17984
rect 7889 17924 7893 17980
rect 7893 17924 7949 17980
rect 7949 17924 7953 17980
rect 7889 17920 7953 17924
rect 7969 17980 8033 17984
rect 7969 17924 7973 17980
rect 7973 17924 8029 17980
rect 8029 17924 8033 17980
rect 7969 17920 8033 17924
rect 14506 17980 14570 17984
rect 14506 17924 14510 17980
rect 14510 17924 14566 17980
rect 14566 17924 14570 17980
rect 14506 17920 14570 17924
rect 14586 17980 14650 17984
rect 14586 17924 14590 17980
rect 14590 17924 14646 17980
rect 14646 17924 14650 17980
rect 14586 17920 14650 17924
rect 14666 17980 14730 17984
rect 14666 17924 14670 17980
rect 14670 17924 14726 17980
rect 14726 17924 14730 17980
rect 14666 17920 14730 17924
rect 14746 17980 14810 17984
rect 14746 17924 14750 17980
rect 14750 17924 14806 17980
rect 14806 17924 14810 17980
rect 14746 17920 14810 17924
rect 4340 17436 4404 17440
rect 4340 17380 4344 17436
rect 4344 17380 4400 17436
rect 4400 17380 4404 17436
rect 4340 17376 4404 17380
rect 4420 17436 4484 17440
rect 4420 17380 4424 17436
rect 4424 17380 4480 17436
rect 4480 17380 4484 17436
rect 4420 17376 4484 17380
rect 4500 17436 4564 17440
rect 4500 17380 4504 17436
rect 4504 17380 4560 17436
rect 4560 17380 4564 17436
rect 4500 17376 4564 17380
rect 4580 17436 4644 17440
rect 4580 17380 4584 17436
rect 4584 17380 4640 17436
rect 4640 17380 4644 17436
rect 4580 17376 4644 17380
rect 11118 17436 11182 17440
rect 11118 17380 11122 17436
rect 11122 17380 11178 17436
rect 11178 17380 11182 17436
rect 11118 17376 11182 17380
rect 11198 17436 11262 17440
rect 11198 17380 11202 17436
rect 11202 17380 11258 17436
rect 11258 17380 11262 17436
rect 11198 17376 11262 17380
rect 11278 17436 11342 17440
rect 11278 17380 11282 17436
rect 11282 17380 11338 17436
rect 11338 17380 11342 17436
rect 11278 17376 11342 17380
rect 11358 17436 11422 17440
rect 11358 17380 11362 17436
rect 11362 17380 11418 17436
rect 11418 17380 11422 17436
rect 11358 17376 11422 17380
rect 17895 17436 17959 17440
rect 17895 17380 17899 17436
rect 17899 17380 17955 17436
rect 17955 17380 17959 17436
rect 17895 17376 17959 17380
rect 17975 17436 18039 17440
rect 17975 17380 17979 17436
rect 17979 17380 18035 17436
rect 18035 17380 18039 17436
rect 17975 17376 18039 17380
rect 18055 17436 18119 17440
rect 18055 17380 18059 17436
rect 18059 17380 18115 17436
rect 18115 17380 18119 17436
rect 18055 17376 18119 17380
rect 18135 17436 18199 17440
rect 18135 17380 18139 17436
rect 18139 17380 18195 17436
rect 18195 17380 18199 17436
rect 18135 17376 18199 17380
rect 7729 16892 7793 16896
rect 7729 16836 7733 16892
rect 7733 16836 7789 16892
rect 7789 16836 7793 16892
rect 7729 16832 7793 16836
rect 7809 16892 7873 16896
rect 7809 16836 7813 16892
rect 7813 16836 7869 16892
rect 7869 16836 7873 16892
rect 7809 16832 7873 16836
rect 7889 16892 7953 16896
rect 7889 16836 7893 16892
rect 7893 16836 7949 16892
rect 7949 16836 7953 16892
rect 7889 16832 7953 16836
rect 7969 16892 8033 16896
rect 7969 16836 7973 16892
rect 7973 16836 8029 16892
rect 8029 16836 8033 16892
rect 7969 16832 8033 16836
rect 14506 16892 14570 16896
rect 14506 16836 14510 16892
rect 14510 16836 14566 16892
rect 14566 16836 14570 16892
rect 14506 16832 14570 16836
rect 14586 16892 14650 16896
rect 14586 16836 14590 16892
rect 14590 16836 14646 16892
rect 14646 16836 14650 16892
rect 14586 16832 14650 16836
rect 14666 16892 14730 16896
rect 14666 16836 14670 16892
rect 14670 16836 14726 16892
rect 14726 16836 14730 16892
rect 14666 16832 14730 16836
rect 14746 16892 14810 16896
rect 14746 16836 14750 16892
rect 14750 16836 14806 16892
rect 14806 16836 14810 16892
rect 14746 16832 14810 16836
rect 4340 16348 4404 16352
rect 4340 16292 4344 16348
rect 4344 16292 4400 16348
rect 4400 16292 4404 16348
rect 4340 16288 4404 16292
rect 4420 16348 4484 16352
rect 4420 16292 4424 16348
rect 4424 16292 4480 16348
rect 4480 16292 4484 16348
rect 4420 16288 4484 16292
rect 4500 16348 4564 16352
rect 4500 16292 4504 16348
rect 4504 16292 4560 16348
rect 4560 16292 4564 16348
rect 4500 16288 4564 16292
rect 4580 16348 4644 16352
rect 4580 16292 4584 16348
rect 4584 16292 4640 16348
rect 4640 16292 4644 16348
rect 4580 16288 4644 16292
rect 11118 16348 11182 16352
rect 11118 16292 11122 16348
rect 11122 16292 11178 16348
rect 11178 16292 11182 16348
rect 11118 16288 11182 16292
rect 11198 16348 11262 16352
rect 11198 16292 11202 16348
rect 11202 16292 11258 16348
rect 11258 16292 11262 16348
rect 11198 16288 11262 16292
rect 11278 16348 11342 16352
rect 11278 16292 11282 16348
rect 11282 16292 11338 16348
rect 11338 16292 11342 16348
rect 11278 16288 11342 16292
rect 11358 16348 11422 16352
rect 11358 16292 11362 16348
rect 11362 16292 11418 16348
rect 11418 16292 11422 16348
rect 11358 16288 11422 16292
rect 17895 16348 17959 16352
rect 17895 16292 17899 16348
rect 17899 16292 17955 16348
rect 17955 16292 17959 16348
rect 17895 16288 17959 16292
rect 17975 16348 18039 16352
rect 17975 16292 17979 16348
rect 17979 16292 18035 16348
rect 18035 16292 18039 16348
rect 17975 16288 18039 16292
rect 18055 16348 18119 16352
rect 18055 16292 18059 16348
rect 18059 16292 18115 16348
rect 18115 16292 18119 16348
rect 18055 16288 18119 16292
rect 18135 16348 18199 16352
rect 18135 16292 18139 16348
rect 18139 16292 18195 16348
rect 18195 16292 18199 16348
rect 18135 16288 18199 16292
rect 7729 15804 7793 15808
rect 7729 15748 7733 15804
rect 7733 15748 7789 15804
rect 7789 15748 7793 15804
rect 7729 15744 7793 15748
rect 7809 15804 7873 15808
rect 7809 15748 7813 15804
rect 7813 15748 7869 15804
rect 7869 15748 7873 15804
rect 7809 15744 7873 15748
rect 7889 15804 7953 15808
rect 7889 15748 7893 15804
rect 7893 15748 7949 15804
rect 7949 15748 7953 15804
rect 7889 15744 7953 15748
rect 7969 15804 8033 15808
rect 7969 15748 7973 15804
rect 7973 15748 8029 15804
rect 8029 15748 8033 15804
rect 7969 15744 8033 15748
rect 14506 15804 14570 15808
rect 14506 15748 14510 15804
rect 14510 15748 14566 15804
rect 14566 15748 14570 15804
rect 14506 15744 14570 15748
rect 14586 15804 14650 15808
rect 14586 15748 14590 15804
rect 14590 15748 14646 15804
rect 14646 15748 14650 15804
rect 14586 15744 14650 15748
rect 14666 15804 14730 15808
rect 14666 15748 14670 15804
rect 14670 15748 14726 15804
rect 14726 15748 14730 15804
rect 14666 15744 14730 15748
rect 14746 15804 14810 15808
rect 14746 15748 14750 15804
rect 14750 15748 14806 15804
rect 14806 15748 14810 15804
rect 14746 15744 14810 15748
rect 4340 15260 4404 15264
rect 4340 15204 4344 15260
rect 4344 15204 4400 15260
rect 4400 15204 4404 15260
rect 4340 15200 4404 15204
rect 4420 15260 4484 15264
rect 4420 15204 4424 15260
rect 4424 15204 4480 15260
rect 4480 15204 4484 15260
rect 4420 15200 4484 15204
rect 4500 15260 4564 15264
rect 4500 15204 4504 15260
rect 4504 15204 4560 15260
rect 4560 15204 4564 15260
rect 4500 15200 4564 15204
rect 4580 15260 4644 15264
rect 4580 15204 4584 15260
rect 4584 15204 4640 15260
rect 4640 15204 4644 15260
rect 4580 15200 4644 15204
rect 11118 15260 11182 15264
rect 11118 15204 11122 15260
rect 11122 15204 11178 15260
rect 11178 15204 11182 15260
rect 11118 15200 11182 15204
rect 11198 15260 11262 15264
rect 11198 15204 11202 15260
rect 11202 15204 11258 15260
rect 11258 15204 11262 15260
rect 11198 15200 11262 15204
rect 11278 15260 11342 15264
rect 11278 15204 11282 15260
rect 11282 15204 11338 15260
rect 11338 15204 11342 15260
rect 11278 15200 11342 15204
rect 11358 15260 11422 15264
rect 11358 15204 11362 15260
rect 11362 15204 11418 15260
rect 11418 15204 11422 15260
rect 11358 15200 11422 15204
rect 17895 15260 17959 15264
rect 17895 15204 17899 15260
rect 17899 15204 17955 15260
rect 17955 15204 17959 15260
rect 17895 15200 17959 15204
rect 17975 15260 18039 15264
rect 17975 15204 17979 15260
rect 17979 15204 18035 15260
rect 18035 15204 18039 15260
rect 17975 15200 18039 15204
rect 18055 15260 18119 15264
rect 18055 15204 18059 15260
rect 18059 15204 18115 15260
rect 18115 15204 18119 15260
rect 18055 15200 18119 15204
rect 18135 15260 18199 15264
rect 18135 15204 18139 15260
rect 18139 15204 18195 15260
rect 18195 15204 18199 15260
rect 18135 15200 18199 15204
rect 7729 14716 7793 14720
rect 7729 14660 7733 14716
rect 7733 14660 7789 14716
rect 7789 14660 7793 14716
rect 7729 14656 7793 14660
rect 7809 14716 7873 14720
rect 7809 14660 7813 14716
rect 7813 14660 7869 14716
rect 7869 14660 7873 14716
rect 7809 14656 7873 14660
rect 7889 14716 7953 14720
rect 7889 14660 7893 14716
rect 7893 14660 7949 14716
rect 7949 14660 7953 14716
rect 7889 14656 7953 14660
rect 7969 14716 8033 14720
rect 7969 14660 7973 14716
rect 7973 14660 8029 14716
rect 8029 14660 8033 14716
rect 7969 14656 8033 14660
rect 14506 14716 14570 14720
rect 14506 14660 14510 14716
rect 14510 14660 14566 14716
rect 14566 14660 14570 14716
rect 14506 14656 14570 14660
rect 14586 14716 14650 14720
rect 14586 14660 14590 14716
rect 14590 14660 14646 14716
rect 14646 14660 14650 14716
rect 14586 14656 14650 14660
rect 14666 14716 14730 14720
rect 14666 14660 14670 14716
rect 14670 14660 14726 14716
rect 14726 14660 14730 14716
rect 14666 14656 14730 14660
rect 14746 14716 14810 14720
rect 14746 14660 14750 14716
rect 14750 14660 14806 14716
rect 14806 14660 14810 14716
rect 14746 14656 14810 14660
rect 4340 14172 4404 14176
rect 4340 14116 4344 14172
rect 4344 14116 4400 14172
rect 4400 14116 4404 14172
rect 4340 14112 4404 14116
rect 4420 14172 4484 14176
rect 4420 14116 4424 14172
rect 4424 14116 4480 14172
rect 4480 14116 4484 14172
rect 4420 14112 4484 14116
rect 4500 14172 4564 14176
rect 4500 14116 4504 14172
rect 4504 14116 4560 14172
rect 4560 14116 4564 14172
rect 4500 14112 4564 14116
rect 4580 14172 4644 14176
rect 4580 14116 4584 14172
rect 4584 14116 4640 14172
rect 4640 14116 4644 14172
rect 4580 14112 4644 14116
rect 11118 14172 11182 14176
rect 11118 14116 11122 14172
rect 11122 14116 11178 14172
rect 11178 14116 11182 14172
rect 11118 14112 11182 14116
rect 11198 14172 11262 14176
rect 11198 14116 11202 14172
rect 11202 14116 11258 14172
rect 11258 14116 11262 14172
rect 11198 14112 11262 14116
rect 11278 14172 11342 14176
rect 11278 14116 11282 14172
rect 11282 14116 11338 14172
rect 11338 14116 11342 14172
rect 11278 14112 11342 14116
rect 11358 14172 11422 14176
rect 11358 14116 11362 14172
rect 11362 14116 11418 14172
rect 11418 14116 11422 14172
rect 11358 14112 11422 14116
rect 17895 14172 17959 14176
rect 17895 14116 17899 14172
rect 17899 14116 17955 14172
rect 17955 14116 17959 14172
rect 17895 14112 17959 14116
rect 17975 14172 18039 14176
rect 17975 14116 17979 14172
rect 17979 14116 18035 14172
rect 18035 14116 18039 14172
rect 17975 14112 18039 14116
rect 18055 14172 18119 14176
rect 18055 14116 18059 14172
rect 18059 14116 18115 14172
rect 18115 14116 18119 14172
rect 18055 14112 18119 14116
rect 18135 14172 18199 14176
rect 18135 14116 18139 14172
rect 18139 14116 18195 14172
rect 18195 14116 18199 14172
rect 18135 14112 18199 14116
rect 7729 13628 7793 13632
rect 7729 13572 7733 13628
rect 7733 13572 7789 13628
rect 7789 13572 7793 13628
rect 7729 13568 7793 13572
rect 7809 13628 7873 13632
rect 7809 13572 7813 13628
rect 7813 13572 7869 13628
rect 7869 13572 7873 13628
rect 7809 13568 7873 13572
rect 7889 13628 7953 13632
rect 7889 13572 7893 13628
rect 7893 13572 7949 13628
rect 7949 13572 7953 13628
rect 7889 13568 7953 13572
rect 7969 13628 8033 13632
rect 7969 13572 7973 13628
rect 7973 13572 8029 13628
rect 8029 13572 8033 13628
rect 7969 13568 8033 13572
rect 14506 13628 14570 13632
rect 14506 13572 14510 13628
rect 14510 13572 14566 13628
rect 14566 13572 14570 13628
rect 14506 13568 14570 13572
rect 14586 13628 14650 13632
rect 14586 13572 14590 13628
rect 14590 13572 14646 13628
rect 14646 13572 14650 13628
rect 14586 13568 14650 13572
rect 14666 13628 14730 13632
rect 14666 13572 14670 13628
rect 14670 13572 14726 13628
rect 14726 13572 14730 13628
rect 14666 13568 14730 13572
rect 14746 13628 14810 13632
rect 14746 13572 14750 13628
rect 14750 13572 14806 13628
rect 14806 13572 14810 13628
rect 14746 13568 14810 13572
rect 4340 13084 4404 13088
rect 4340 13028 4344 13084
rect 4344 13028 4400 13084
rect 4400 13028 4404 13084
rect 4340 13024 4404 13028
rect 4420 13084 4484 13088
rect 4420 13028 4424 13084
rect 4424 13028 4480 13084
rect 4480 13028 4484 13084
rect 4420 13024 4484 13028
rect 4500 13084 4564 13088
rect 4500 13028 4504 13084
rect 4504 13028 4560 13084
rect 4560 13028 4564 13084
rect 4500 13024 4564 13028
rect 4580 13084 4644 13088
rect 4580 13028 4584 13084
rect 4584 13028 4640 13084
rect 4640 13028 4644 13084
rect 4580 13024 4644 13028
rect 11118 13084 11182 13088
rect 11118 13028 11122 13084
rect 11122 13028 11178 13084
rect 11178 13028 11182 13084
rect 11118 13024 11182 13028
rect 11198 13084 11262 13088
rect 11198 13028 11202 13084
rect 11202 13028 11258 13084
rect 11258 13028 11262 13084
rect 11198 13024 11262 13028
rect 11278 13084 11342 13088
rect 11278 13028 11282 13084
rect 11282 13028 11338 13084
rect 11338 13028 11342 13084
rect 11278 13024 11342 13028
rect 11358 13084 11422 13088
rect 11358 13028 11362 13084
rect 11362 13028 11418 13084
rect 11418 13028 11422 13084
rect 11358 13024 11422 13028
rect 17895 13084 17959 13088
rect 17895 13028 17899 13084
rect 17899 13028 17955 13084
rect 17955 13028 17959 13084
rect 17895 13024 17959 13028
rect 17975 13084 18039 13088
rect 17975 13028 17979 13084
rect 17979 13028 18035 13084
rect 18035 13028 18039 13084
rect 17975 13024 18039 13028
rect 18055 13084 18119 13088
rect 18055 13028 18059 13084
rect 18059 13028 18115 13084
rect 18115 13028 18119 13084
rect 18055 13024 18119 13028
rect 18135 13084 18199 13088
rect 18135 13028 18139 13084
rect 18139 13028 18195 13084
rect 18195 13028 18199 13084
rect 18135 13024 18199 13028
rect 7729 12540 7793 12544
rect 7729 12484 7733 12540
rect 7733 12484 7789 12540
rect 7789 12484 7793 12540
rect 7729 12480 7793 12484
rect 7809 12540 7873 12544
rect 7809 12484 7813 12540
rect 7813 12484 7869 12540
rect 7869 12484 7873 12540
rect 7809 12480 7873 12484
rect 7889 12540 7953 12544
rect 7889 12484 7893 12540
rect 7893 12484 7949 12540
rect 7949 12484 7953 12540
rect 7889 12480 7953 12484
rect 7969 12540 8033 12544
rect 7969 12484 7973 12540
rect 7973 12484 8029 12540
rect 8029 12484 8033 12540
rect 7969 12480 8033 12484
rect 14506 12540 14570 12544
rect 14506 12484 14510 12540
rect 14510 12484 14566 12540
rect 14566 12484 14570 12540
rect 14506 12480 14570 12484
rect 14586 12540 14650 12544
rect 14586 12484 14590 12540
rect 14590 12484 14646 12540
rect 14646 12484 14650 12540
rect 14586 12480 14650 12484
rect 14666 12540 14730 12544
rect 14666 12484 14670 12540
rect 14670 12484 14726 12540
rect 14726 12484 14730 12540
rect 14666 12480 14730 12484
rect 14746 12540 14810 12544
rect 14746 12484 14750 12540
rect 14750 12484 14806 12540
rect 14806 12484 14810 12540
rect 14746 12480 14810 12484
rect 4340 11996 4404 12000
rect 4340 11940 4344 11996
rect 4344 11940 4400 11996
rect 4400 11940 4404 11996
rect 4340 11936 4404 11940
rect 4420 11996 4484 12000
rect 4420 11940 4424 11996
rect 4424 11940 4480 11996
rect 4480 11940 4484 11996
rect 4420 11936 4484 11940
rect 4500 11996 4564 12000
rect 4500 11940 4504 11996
rect 4504 11940 4560 11996
rect 4560 11940 4564 11996
rect 4500 11936 4564 11940
rect 4580 11996 4644 12000
rect 4580 11940 4584 11996
rect 4584 11940 4640 11996
rect 4640 11940 4644 11996
rect 4580 11936 4644 11940
rect 11118 11996 11182 12000
rect 11118 11940 11122 11996
rect 11122 11940 11178 11996
rect 11178 11940 11182 11996
rect 11118 11936 11182 11940
rect 11198 11996 11262 12000
rect 11198 11940 11202 11996
rect 11202 11940 11258 11996
rect 11258 11940 11262 11996
rect 11198 11936 11262 11940
rect 11278 11996 11342 12000
rect 11278 11940 11282 11996
rect 11282 11940 11338 11996
rect 11338 11940 11342 11996
rect 11278 11936 11342 11940
rect 11358 11996 11422 12000
rect 11358 11940 11362 11996
rect 11362 11940 11418 11996
rect 11418 11940 11422 11996
rect 11358 11936 11422 11940
rect 17895 11996 17959 12000
rect 17895 11940 17899 11996
rect 17899 11940 17955 11996
rect 17955 11940 17959 11996
rect 17895 11936 17959 11940
rect 17975 11996 18039 12000
rect 17975 11940 17979 11996
rect 17979 11940 18035 11996
rect 18035 11940 18039 11996
rect 17975 11936 18039 11940
rect 18055 11996 18119 12000
rect 18055 11940 18059 11996
rect 18059 11940 18115 11996
rect 18115 11940 18119 11996
rect 18055 11936 18119 11940
rect 18135 11996 18199 12000
rect 18135 11940 18139 11996
rect 18139 11940 18195 11996
rect 18195 11940 18199 11996
rect 18135 11936 18199 11940
rect 7729 11452 7793 11456
rect 7729 11396 7733 11452
rect 7733 11396 7789 11452
rect 7789 11396 7793 11452
rect 7729 11392 7793 11396
rect 7809 11452 7873 11456
rect 7809 11396 7813 11452
rect 7813 11396 7869 11452
rect 7869 11396 7873 11452
rect 7809 11392 7873 11396
rect 7889 11452 7953 11456
rect 7889 11396 7893 11452
rect 7893 11396 7949 11452
rect 7949 11396 7953 11452
rect 7889 11392 7953 11396
rect 7969 11452 8033 11456
rect 7969 11396 7973 11452
rect 7973 11396 8029 11452
rect 8029 11396 8033 11452
rect 7969 11392 8033 11396
rect 14506 11452 14570 11456
rect 14506 11396 14510 11452
rect 14510 11396 14566 11452
rect 14566 11396 14570 11452
rect 14506 11392 14570 11396
rect 14586 11452 14650 11456
rect 14586 11396 14590 11452
rect 14590 11396 14646 11452
rect 14646 11396 14650 11452
rect 14586 11392 14650 11396
rect 14666 11452 14730 11456
rect 14666 11396 14670 11452
rect 14670 11396 14726 11452
rect 14726 11396 14730 11452
rect 14666 11392 14730 11396
rect 14746 11452 14810 11456
rect 14746 11396 14750 11452
rect 14750 11396 14806 11452
rect 14806 11396 14810 11452
rect 14746 11392 14810 11396
rect 4340 10908 4404 10912
rect 4340 10852 4344 10908
rect 4344 10852 4400 10908
rect 4400 10852 4404 10908
rect 4340 10848 4404 10852
rect 4420 10908 4484 10912
rect 4420 10852 4424 10908
rect 4424 10852 4480 10908
rect 4480 10852 4484 10908
rect 4420 10848 4484 10852
rect 4500 10908 4564 10912
rect 4500 10852 4504 10908
rect 4504 10852 4560 10908
rect 4560 10852 4564 10908
rect 4500 10848 4564 10852
rect 4580 10908 4644 10912
rect 4580 10852 4584 10908
rect 4584 10852 4640 10908
rect 4640 10852 4644 10908
rect 4580 10848 4644 10852
rect 11118 10908 11182 10912
rect 11118 10852 11122 10908
rect 11122 10852 11178 10908
rect 11178 10852 11182 10908
rect 11118 10848 11182 10852
rect 11198 10908 11262 10912
rect 11198 10852 11202 10908
rect 11202 10852 11258 10908
rect 11258 10852 11262 10908
rect 11198 10848 11262 10852
rect 11278 10908 11342 10912
rect 11278 10852 11282 10908
rect 11282 10852 11338 10908
rect 11338 10852 11342 10908
rect 11278 10848 11342 10852
rect 11358 10908 11422 10912
rect 11358 10852 11362 10908
rect 11362 10852 11418 10908
rect 11418 10852 11422 10908
rect 11358 10848 11422 10852
rect 17895 10908 17959 10912
rect 17895 10852 17899 10908
rect 17899 10852 17955 10908
rect 17955 10852 17959 10908
rect 17895 10848 17959 10852
rect 17975 10908 18039 10912
rect 17975 10852 17979 10908
rect 17979 10852 18035 10908
rect 18035 10852 18039 10908
rect 17975 10848 18039 10852
rect 18055 10908 18119 10912
rect 18055 10852 18059 10908
rect 18059 10852 18115 10908
rect 18115 10852 18119 10908
rect 18055 10848 18119 10852
rect 18135 10908 18199 10912
rect 18135 10852 18139 10908
rect 18139 10852 18195 10908
rect 18195 10852 18199 10908
rect 18135 10848 18199 10852
rect 7729 10364 7793 10368
rect 7729 10308 7733 10364
rect 7733 10308 7789 10364
rect 7789 10308 7793 10364
rect 7729 10304 7793 10308
rect 7809 10364 7873 10368
rect 7809 10308 7813 10364
rect 7813 10308 7869 10364
rect 7869 10308 7873 10364
rect 7809 10304 7873 10308
rect 7889 10364 7953 10368
rect 7889 10308 7893 10364
rect 7893 10308 7949 10364
rect 7949 10308 7953 10364
rect 7889 10304 7953 10308
rect 7969 10364 8033 10368
rect 7969 10308 7973 10364
rect 7973 10308 8029 10364
rect 8029 10308 8033 10364
rect 7969 10304 8033 10308
rect 14506 10364 14570 10368
rect 14506 10308 14510 10364
rect 14510 10308 14566 10364
rect 14566 10308 14570 10364
rect 14506 10304 14570 10308
rect 14586 10364 14650 10368
rect 14586 10308 14590 10364
rect 14590 10308 14646 10364
rect 14646 10308 14650 10364
rect 14586 10304 14650 10308
rect 14666 10364 14730 10368
rect 14666 10308 14670 10364
rect 14670 10308 14726 10364
rect 14726 10308 14730 10364
rect 14666 10304 14730 10308
rect 14746 10364 14810 10368
rect 14746 10308 14750 10364
rect 14750 10308 14806 10364
rect 14806 10308 14810 10364
rect 14746 10304 14810 10308
rect 4340 9820 4404 9824
rect 4340 9764 4344 9820
rect 4344 9764 4400 9820
rect 4400 9764 4404 9820
rect 4340 9760 4404 9764
rect 4420 9820 4484 9824
rect 4420 9764 4424 9820
rect 4424 9764 4480 9820
rect 4480 9764 4484 9820
rect 4420 9760 4484 9764
rect 4500 9820 4564 9824
rect 4500 9764 4504 9820
rect 4504 9764 4560 9820
rect 4560 9764 4564 9820
rect 4500 9760 4564 9764
rect 4580 9820 4644 9824
rect 4580 9764 4584 9820
rect 4584 9764 4640 9820
rect 4640 9764 4644 9820
rect 4580 9760 4644 9764
rect 11118 9820 11182 9824
rect 11118 9764 11122 9820
rect 11122 9764 11178 9820
rect 11178 9764 11182 9820
rect 11118 9760 11182 9764
rect 11198 9820 11262 9824
rect 11198 9764 11202 9820
rect 11202 9764 11258 9820
rect 11258 9764 11262 9820
rect 11198 9760 11262 9764
rect 11278 9820 11342 9824
rect 11278 9764 11282 9820
rect 11282 9764 11338 9820
rect 11338 9764 11342 9820
rect 11278 9760 11342 9764
rect 11358 9820 11422 9824
rect 11358 9764 11362 9820
rect 11362 9764 11418 9820
rect 11418 9764 11422 9820
rect 11358 9760 11422 9764
rect 17895 9820 17959 9824
rect 17895 9764 17899 9820
rect 17899 9764 17955 9820
rect 17955 9764 17959 9820
rect 17895 9760 17959 9764
rect 17975 9820 18039 9824
rect 17975 9764 17979 9820
rect 17979 9764 18035 9820
rect 18035 9764 18039 9820
rect 17975 9760 18039 9764
rect 18055 9820 18119 9824
rect 18055 9764 18059 9820
rect 18059 9764 18115 9820
rect 18115 9764 18119 9820
rect 18055 9760 18119 9764
rect 18135 9820 18199 9824
rect 18135 9764 18139 9820
rect 18139 9764 18195 9820
rect 18195 9764 18199 9820
rect 18135 9760 18199 9764
rect 7729 9276 7793 9280
rect 7729 9220 7733 9276
rect 7733 9220 7789 9276
rect 7789 9220 7793 9276
rect 7729 9216 7793 9220
rect 7809 9276 7873 9280
rect 7809 9220 7813 9276
rect 7813 9220 7869 9276
rect 7869 9220 7873 9276
rect 7809 9216 7873 9220
rect 7889 9276 7953 9280
rect 7889 9220 7893 9276
rect 7893 9220 7949 9276
rect 7949 9220 7953 9276
rect 7889 9216 7953 9220
rect 7969 9276 8033 9280
rect 7969 9220 7973 9276
rect 7973 9220 8029 9276
rect 8029 9220 8033 9276
rect 7969 9216 8033 9220
rect 14506 9276 14570 9280
rect 14506 9220 14510 9276
rect 14510 9220 14566 9276
rect 14566 9220 14570 9276
rect 14506 9216 14570 9220
rect 14586 9276 14650 9280
rect 14586 9220 14590 9276
rect 14590 9220 14646 9276
rect 14646 9220 14650 9276
rect 14586 9216 14650 9220
rect 14666 9276 14730 9280
rect 14666 9220 14670 9276
rect 14670 9220 14726 9276
rect 14726 9220 14730 9276
rect 14666 9216 14730 9220
rect 14746 9276 14810 9280
rect 14746 9220 14750 9276
rect 14750 9220 14806 9276
rect 14806 9220 14810 9276
rect 14746 9216 14810 9220
rect 4340 8732 4404 8736
rect 4340 8676 4344 8732
rect 4344 8676 4400 8732
rect 4400 8676 4404 8732
rect 4340 8672 4404 8676
rect 4420 8732 4484 8736
rect 4420 8676 4424 8732
rect 4424 8676 4480 8732
rect 4480 8676 4484 8732
rect 4420 8672 4484 8676
rect 4500 8732 4564 8736
rect 4500 8676 4504 8732
rect 4504 8676 4560 8732
rect 4560 8676 4564 8732
rect 4500 8672 4564 8676
rect 4580 8732 4644 8736
rect 4580 8676 4584 8732
rect 4584 8676 4640 8732
rect 4640 8676 4644 8732
rect 4580 8672 4644 8676
rect 11118 8732 11182 8736
rect 11118 8676 11122 8732
rect 11122 8676 11178 8732
rect 11178 8676 11182 8732
rect 11118 8672 11182 8676
rect 11198 8732 11262 8736
rect 11198 8676 11202 8732
rect 11202 8676 11258 8732
rect 11258 8676 11262 8732
rect 11198 8672 11262 8676
rect 11278 8732 11342 8736
rect 11278 8676 11282 8732
rect 11282 8676 11338 8732
rect 11338 8676 11342 8732
rect 11278 8672 11342 8676
rect 11358 8732 11422 8736
rect 11358 8676 11362 8732
rect 11362 8676 11418 8732
rect 11418 8676 11422 8732
rect 11358 8672 11422 8676
rect 17895 8732 17959 8736
rect 17895 8676 17899 8732
rect 17899 8676 17955 8732
rect 17955 8676 17959 8732
rect 17895 8672 17959 8676
rect 17975 8732 18039 8736
rect 17975 8676 17979 8732
rect 17979 8676 18035 8732
rect 18035 8676 18039 8732
rect 17975 8672 18039 8676
rect 18055 8732 18119 8736
rect 18055 8676 18059 8732
rect 18059 8676 18115 8732
rect 18115 8676 18119 8732
rect 18055 8672 18119 8676
rect 18135 8732 18199 8736
rect 18135 8676 18139 8732
rect 18139 8676 18195 8732
rect 18195 8676 18199 8732
rect 18135 8672 18199 8676
rect 7729 8188 7793 8192
rect 7729 8132 7733 8188
rect 7733 8132 7789 8188
rect 7789 8132 7793 8188
rect 7729 8128 7793 8132
rect 7809 8188 7873 8192
rect 7809 8132 7813 8188
rect 7813 8132 7869 8188
rect 7869 8132 7873 8188
rect 7809 8128 7873 8132
rect 7889 8188 7953 8192
rect 7889 8132 7893 8188
rect 7893 8132 7949 8188
rect 7949 8132 7953 8188
rect 7889 8128 7953 8132
rect 7969 8188 8033 8192
rect 7969 8132 7973 8188
rect 7973 8132 8029 8188
rect 8029 8132 8033 8188
rect 7969 8128 8033 8132
rect 14506 8188 14570 8192
rect 14506 8132 14510 8188
rect 14510 8132 14566 8188
rect 14566 8132 14570 8188
rect 14506 8128 14570 8132
rect 14586 8188 14650 8192
rect 14586 8132 14590 8188
rect 14590 8132 14646 8188
rect 14646 8132 14650 8188
rect 14586 8128 14650 8132
rect 14666 8188 14730 8192
rect 14666 8132 14670 8188
rect 14670 8132 14726 8188
rect 14726 8132 14730 8188
rect 14666 8128 14730 8132
rect 14746 8188 14810 8192
rect 14746 8132 14750 8188
rect 14750 8132 14806 8188
rect 14806 8132 14810 8188
rect 14746 8128 14810 8132
rect 4340 7644 4404 7648
rect 4340 7588 4344 7644
rect 4344 7588 4400 7644
rect 4400 7588 4404 7644
rect 4340 7584 4404 7588
rect 4420 7644 4484 7648
rect 4420 7588 4424 7644
rect 4424 7588 4480 7644
rect 4480 7588 4484 7644
rect 4420 7584 4484 7588
rect 4500 7644 4564 7648
rect 4500 7588 4504 7644
rect 4504 7588 4560 7644
rect 4560 7588 4564 7644
rect 4500 7584 4564 7588
rect 4580 7644 4644 7648
rect 4580 7588 4584 7644
rect 4584 7588 4640 7644
rect 4640 7588 4644 7644
rect 4580 7584 4644 7588
rect 11118 7644 11182 7648
rect 11118 7588 11122 7644
rect 11122 7588 11178 7644
rect 11178 7588 11182 7644
rect 11118 7584 11182 7588
rect 11198 7644 11262 7648
rect 11198 7588 11202 7644
rect 11202 7588 11258 7644
rect 11258 7588 11262 7644
rect 11198 7584 11262 7588
rect 11278 7644 11342 7648
rect 11278 7588 11282 7644
rect 11282 7588 11338 7644
rect 11338 7588 11342 7644
rect 11278 7584 11342 7588
rect 11358 7644 11422 7648
rect 11358 7588 11362 7644
rect 11362 7588 11418 7644
rect 11418 7588 11422 7644
rect 11358 7584 11422 7588
rect 17895 7644 17959 7648
rect 17895 7588 17899 7644
rect 17899 7588 17955 7644
rect 17955 7588 17959 7644
rect 17895 7584 17959 7588
rect 17975 7644 18039 7648
rect 17975 7588 17979 7644
rect 17979 7588 18035 7644
rect 18035 7588 18039 7644
rect 17975 7584 18039 7588
rect 18055 7644 18119 7648
rect 18055 7588 18059 7644
rect 18059 7588 18115 7644
rect 18115 7588 18119 7644
rect 18055 7584 18119 7588
rect 18135 7644 18199 7648
rect 18135 7588 18139 7644
rect 18139 7588 18195 7644
rect 18195 7588 18199 7644
rect 18135 7584 18199 7588
rect 7729 7100 7793 7104
rect 7729 7044 7733 7100
rect 7733 7044 7789 7100
rect 7789 7044 7793 7100
rect 7729 7040 7793 7044
rect 7809 7100 7873 7104
rect 7809 7044 7813 7100
rect 7813 7044 7869 7100
rect 7869 7044 7873 7100
rect 7809 7040 7873 7044
rect 7889 7100 7953 7104
rect 7889 7044 7893 7100
rect 7893 7044 7949 7100
rect 7949 7044 7953 7100
rect 7889 7040 7953 7044
rect 7969 7100 8033 7104
rect 7969 7044 7973 7100
rect 7973 7044 8029 7100
rect 8029 7044 8033 7100
rect 7969 7040 8033 7044
rect 14506 7100 14570 7104
rect 14506 7044 14510 7100
rect 14510 7044 14566 7100
rect 14566 7044 14570 7100
rect 14506 7040 14570 7044
rect 14586 7100 14650 7104
rect 14586 7044 14590 7100
rect 14590 7044 14646 7100
rect 14646 7044 14650 7100
rect 14586 7040 14650 7044
rect 14666 7100 14730 7104
rect 14666 7044 14670 7100
rect 14670 7044 14726 7100
rect 14726 7044 14730 7100
rect 14666 7040 14730 7044
rect 14746 7100 14810 7104
rect 14746 7044 14750 7100
rect 14750 7044 14806 7100
rect 14806 7044 14810 7100
rect 14746 7040 14810 7044
rect 4340 6556 4404 6560
rect 4340 6500 4344 6556
rect 4344 6500 4400 6556
rect 4400 6500 4404 6556
rect 4340 6496 4404 6500
rect 4420 6556 4484 6560
rect 4420 6500 4424 6556
rect 4424 6500 4480 6556
rect 4480 6500 4484 6556
rect 4420 6496 4484 6500
rect 4500 6556 4564 6560
rect 4500 6500 4504 6556
rect 4504 6500 4560 6556
rect 4560 6500 4564 6556
rect 4500 6496 4564 6500
rect 4580 6556 4644 6560
rect 4580 6500 4584 6556
rect 4584 6500 4640 6556
rect 4640 6500 4644 6556
rect 4580 6496 4644 6500
rect 11118 6556 11182 6560
rect 11118 6500 11122 6556
rect 11122 6500 11178 6556
rect 11178 6500 11182 6556
rect 11118 6496 11182 6500
rect 11198 6556 11262 6560
rect 11198 6500 11202 6556
rect 11202 6500 11258 6556
rect 11258 6500 11262 6556
rect 11198 6496 11262 6500
rect 11278 6556 11342 6560
rect 11278 6500 11282 6556
rect 11282 6500 11338 6556
rect 11338 6500 11342 6556
rect 11278 6496 11342 6500
rect 11358 6556 11422 6560
rect 11358 6500 11362 6556
rect 11362 6500 11418 6556
rect 11418 6500 11422 6556
rect 11358 6496 11422 6500
rect 17895 6556 17959 6560
rect 17895 6500 17899 6556
rect 17899 6500 17955 6556
rect 17955 6500 17959 6556
rect 17895 6496 17959 6500
rect 17975 6556 18039 6560
rect 17975 6500 17979 6556
rect 17979 6500 18035 6556
rect 18035 6500 18039 6556
rect 17975 6496 18039 6500
rect 18055 6556 18119 6560
rect 18055 6500 18059 6556
rect 18059 6500 18115 6556
rect 18115 6500 18119 6556
rect 18055 6496 18119 6500
rect 18135 6556 18199 6560
rect 18135 6500 18139 6556
rect 18139 6500 18195 6556
rect 18195 6500 18199 6556
rect 18135 6496 18199 6500
rect 7729 6012 7793 6016
rect 7729 5956 7733 6012
rect 7733 5956 7789 6012
rect 7789 5956 7793 6012
rect 7729 5952 7793 5956
rect 7809 6012 7873 6016
rect 7809 5956 7813 6012
rect 7813 5956 7869 6012
rect 7869 5956 7873 6012
rect 7809 5952 7873 5956
rect 7889 6012 7953 6016
rect 7889 5956 7893 6012
rect 7893 5956 7949 6012
rect 7949 5956 7953 6012
rect 7889 5952 7953 5956
rect 7969 6012 8033 6016
rect 7969 5956 7973 6012
rect 7973 5956 8029 6012
rect 8029 5956 8033 6012
rect 7969 5952 8033 5956
rect 14506 6012 14570 6016
rect 14506 5956 14510 6012
rect 14510 5956 14566 6012
rect 14566 5956 14570 6012
rect 14506 5952 14570 5956
rect 14586 6012 14650 6016
rect 14586 5956 14590 6012
rect 14590 5956 14646 6012
rect 14646 5956 14650 6012
rect 14586 5952 14650 5956
rect 14666 6012 14730 6016
rect 14666 5956 14670 6012
rect 14670 5956 14726 6012
rect 14726 5956 14730 6012
rect 14666 5952 14730 5956
rect 14746 6012 14810 6016
rect 14746 5956 14750 6012
rect 14750 5956 14806 6012
rect 14806 5956 14810 6012
rect 14746 5952 14810 5956
rect 4340 5468 4404 5472
rect 4340 5412 4344 5468
rect 4344 5412 4400 5468
rect 4400 5412 4404 5468
rect 4340 5408 4404 5412
rect 4420 5468 4484 5472
rect 4420 5412 4424 5468
rect 4424 5412 4480 5468
rect 4480 5412 4484 5468
rect 4420 5408 4484 5412
rect 4500 5468 4564 5472
rect 4500 5412 4504 5468
rect 4504 5412 4560 5468
rect 4560 5412 4564 5468
rect 4500 5408 4564 5412
rect 4580 5468 4644 5472
rect 4580 5412 4584 5468
rect 4584 5412 4640 5468
rect 4640 5412 4644 5468
rect 4580 5408 4644 5412
rect 11118 5468 11182 5472
rect 11118 5412 11122 5468
rect 11122 5412 11178 5468
rect 11178 5412 11182 5468
rect 11118 5408 11182 5412
rect 11198 5468 11262 5472
rect 11198 5412 11202 5468
rect 11202 5412 11258 5468
rect 11258 5412 11262 5468
rect 11198 5408 11262 5412
rect 11278 5468 11342 5472
rect 11278 5412 11282 5468
rect 11282 5412 11338 5468
rect 11338 5412 11342 5468
rect 11278 5408 11342 5412
rect 11358 5468 11422 5472
rect 11358 5412 11362 5468
rect 11362 5412 11418 5468
rect 11418 5412 11422 5468
rect 11358 5408 11422 5412
rect 17895 5468 17959 5472
rect 17895 5412 17899 5468
rect 17899 5412 17955 5468
rect 17955 5412 17959 5468
rect 17895 5408 17959 5412
rect 17975 5468 18039 5472
rect 17975 5412 17979 5468
rect 17979 5412 18035 5468
rect 18035 5412 18039 5468
rect 17975 5408 18039 5412
rect 18055 5468 18119 5472
rect 18055 5412 18059 5468
rect 18059 5412 18115 5468
rect 18115 5412 18119 5468
rect 18055 5408 18119 5412
rect 18135 5468 18199 5472
rect 18135 5412 18139 5468
rect 18139 5412 18195 5468
rect 18195 5412 18199 5468
rect 18135 5408 18199 5412
rect 7729 4924 7793 4928
rect 7729 4868 7733 4924
rect 7733 4868 7789 4924
rect 7789 4868 7793 4924
rect 7729 4864 7793 4868
rect 7809 4924 7873 4928
rect 7809 4868 7813 4924
rect 7813 4868 7869 4924
rect 7869 4868 7873 4924
rect 7809 4864 7873 4868
rect 7889 4924 7953 4928
rect 7889 4868 7893 4924
rect 7893 4868 7949 4924
rect 7949 4868 7953 4924
rect 7889 4864 7953 4868
rect 7969 4924 8033 4928
rect 7969 4868 7973 4924
rect 7973 4868 8029 4924
rect 8029 4868 8033 4924
rect 7969 4864 8033 4868
rect 14506 4924 14570 4928
rect 14506 4868 14510 4924
rect 14510 4868 14566 4924
rect 14566 4868 14570 4924
rect 14506 4864 14570 4868
rect 14586 4924 14650 4928
rect 14586 4868 14590 4924
rect 14590 4868 14646 4924
rect 14646 4868 14650 4924
rect 14586 4864 14650 4868
rect 14666 4924 14730 4928
rect 14666 4868 14670 4924
rect 14670 4868 14726 4924
rect 14726 4868 14730 4924
rect 14666 4864 14730 4868
rect 14746 4924 14810 4928
rect 14746 4868 14750 4924
rect 14750 4868 14806 4924
rect 14806 4868 14810 4924
rect 14746 4864 14810 4868
rect 4340 4380 4404 4384
rect 4340 4324 4344 4380
rect 4344 4324 4400 4380
rect 4400 4324 4404 4380
rect 4340 4320 4404 4324
rect 4420 4380 4484 4384
rect 4420 4324 4424 4380
rect 4424 4324 4480 4380
rect 4480 4324 4484 4380
rect 4420 4320 4484 4324
rect 4500 4380 4564 4384
rect 4500 4324 4504 4380
rect 4504 4324 4560 4380
rect 4560 4324 4564 4380
rect 4500 4320 4564 4324
rect 4580 4380 4644 4384
rect 4580 4324 4584 4380
rect 4584 4324 4640 4380
rect 4640 4324 4644 4380
rect 4580 4320 4644 4324
rect 11118 4380 11182 4384
rect 11118 4324 11122 4380
rect 11122 4324 11178 4380
rect 11178 4324 11182 4380
rect 11118 4320 11182 4324
rect 11198 4380 11262 4384
rect 11198 4324 11202 4380
rect 11202 4324 11258 4380
rect 11258 4324 11262 4380
rect 11198 4320 11262 4324
rect 11278 4380 11342 4384
rect 11278 4324 11282 4380
rect 11282 4324 11338 4380
rect 11338 4324 11342 4380
rect 11278 4320 11342 4324
rect 11358 4380 11422 4384
rect 11358 4324 11362 4380
rect 11362 4324 11418 4380
rect 11418 4324 11422 4380
rect 11358 4320 11422 4324
rect 17895 4380 17959 4384
rect 17895 4324 17899 4380
rect 17899 4324 17955 4380
rect 17955 4324 17959 4380
rect 17895 4320 17959 4324
rect 17975 4380 18039 4384
rect 17975 4324 17979 4380
rect 17979 4324 18035 4380
rect 18035 4324 18039 4380
rect 17975 4320 18039 4324
rect 18055 4380 18119 4384
rect 18055 4324 18059 4380
rect 18059 4324 18115 4380
rect 18115 4324 18119 4380
rect 18055 4320 18119 4324
rect 18135 4380 18199 4384
rect 18135 4324 18139 4380
rect 18139 4324 18195 4380
rect 18195 4324 18199 4380
rect 18135 4320 18199 4324
rect 7729 3836 7793 3840
rect 7729 3780 7733 3836
rect 7733 3780 7789 3836
rect 7789 3780 7793 3836
rect 7729 3776 7793 3780
rect 7809 3836 7873 3840
rect 7809 3780 7813 3836
rect 7813 3780 7869 3836
rect 7869 3780 7873 3836
rect 7809 3776 7873 3780
rect 7889 3836 7953 3840
rect 7889 3780 7893 3836
rect 7893 3780 7949 3836
rect 7949 3780 7953 3836
rect 7889 3776 7953 3780
rect 7969 3836 8033 3840
rect 7969 3780 7973 3836
rect 7973 3780 8029 3836
rect 8029 3780 8033 3836
rect 7969 3776 8033 3780
rect 14506 3836 14570 3840
rect 14506 3780 14510 3836
rect 14510 3780 14566 3836
rect 14566 3780 14570 3836
rect 14506 3776 14570 3780
rect 14586 3836 14650 3840
rect 14586 3780 14590 3836
rect 14590 3780 14646 3836
rect 14646 3780 14650 3836
rect 14586 3776 14650 3780
rect 14666 3836 14730 3840
rect 14666 3780 14670 3836
rect 14670 3780 14726 3836
rect 14726 3780 14730 3836
rect 14666 3776 14730 3780
rect 14746 3836 14810 3840
rect 14746 3780 14750 3836
rect 14750 3780 14806 3836
rect 14806 3780 14810 3836
rect 14746 3776 14810 3780
rect 4340 3292 4404 3296
rect 4340 3236 4344 3292
rect 4344 3236 4400 3292
rect 4400 3236 4404 3292
rect 4340 3232 4404 3236
rect 4420 3292 4484 3296
rect 4420 3236 4424 3292
rect 4424 3236 4480 3292
rect 4480 3236 4484 3292
rect 4420 3232 4484 3236
rect 4500 3292 4564 3296
rect 4500 3236 4504 3292
rect 4504 3236 4560 3292
rect 4560 3236 4564 3292
rect 4500 3232 4564 3236
rect 4580 3292 4644 3296
rect 4580 3236 4584 3292
rect 4584 3236 4640 3292
rect 4640 3236 4644 3292
rect 4580 3232 4644 3236
rect 11118 3292 11182 3296
rect 11118 3236 11122 3292
rect 11122 3236 11178 3292
rect 11178 3236 11182 3292
rect 11118 3232 11182 3236
rect 11198 3292 11262 3296
rect 11198 3236 11202 3292
rect 11202 3236 11258 3292
rect 11258 3236 11262 3292
rect 11198 3232 11262 3236
rect 11278 3292 11342 3296
rect 11278 3236 11282 3292
rect 11282 3236 11338 3292
rect 11338 3236 11342 3292
rect 11278 3232 11342 3236
rect 11358 3292 11422 3296
rect 11358 3236 11362 3292
rect 11362 3236 11418 3292
rect 11418 3236 11422 3292
rect 11358 3232 11422 3236
rect 17895 3292 17959 3296
rect 17895 3236 17899 3292
rect 17899 3236 17955 3292
rect 17955 3236 17959 3292
rect 17895 3232 17959 3236
rect 17975 3292 18039 3296
rect 17975 3236 17979 3292
rect 17979 3236 18035 3292
rect 18035 3236 18039 3292
rect 17975 3232 18039 3236
rect 18055 3292 18119 3296
rect 18055 3236 18059 3292
rect 18059 3236 18115 3292
rect 18115 3236 18119 3292
rect 18055 3232 18119 3236
rect 18135 3292 18199 3296
rect 18135 3236 18139 3292
rect 18139 3236 18195 3292
rect 18195 3236 18199 3292
rect 18135 3232 18199 3236
rect 7729 2748 7793 2752
rect 7729 2692 7733 2748
rect 7733 2692 7789 2748
rect 7789 2692 7793 2748
rect 7729 2688 7793 2692
rect 7809 2748 7873 2752
rect 7809 2692 7813 2748
rect 7813 2692 7869 2748
rect 7869 2692 7873 2748
rect 7809 2688 7873 2692
rect 7889 2748 7953 2752
rect 7889 2692 7893 2748
rect 7893 2692 7949 2748
rect 7949 2692 7953 2748
rect 7889 2688 7953 2692
rect 7969 2748 8033 2752
rect 7969 2692 7973 2748
rect 7973 2692 8029 2748
rect 8029 2692 8033 2748
rect 7969 2688 8033 2692
rect 14506 2748 14570 2752
rect 14506 2692 14510 2748
rect 14510 2692 14566 2748
rect 14566 2692 14570 2748
rect 14506 2688 14570 2692
rect 14586 2748 14650 2752
rect 14586 2692 14590 2748
rect 14590 2692 14646 2748
rect 14646 2692 14650 2748
rect 14586 2688 14650 2692
rect 14666 2748 14730 2752
rect 14666 2692 14670 2748
rect 14670 2692 14726 2748
rect 14726 2692 14730 2748
rect 14666 2688 14730 2692
rect 14746 2748 14810 2752
rect 14746 2692 14750 2748
rect 14750 2692 14806 2748
rect 14806 2692 14810 2748
rect 14746 2688 14810 2692
rect 4340 2204 4404 2208
rect 4340 2148 4344 2204
rect 4344 2148 4400 2204
rect 4400 2148 4404 2204
rect 4340 2144 4404 2148
rect 4420 2204 4484 2208
rect 4420 2148 4424 2204
rect 4424 2148 4480 2204
rect 4480 2148 4484 2204
rect 4420 2144 4484 2148
rect 4500 2204 4564 2208
rect 4500 2148 4504 2204
rect 4504 2148 4560 2204
rect 4560 2148 4564 2204
rect 4500 2144 4564 2148
rect 4580 2204 4644 2208
rect 4580 2148 4584 2204
rect 4584 2148 4640 2204
rect 4640 2148 4644 2204
rect 4580 2144 4644 2148
rect 11118 2204 11182 2208
rect 11118 2148 11122 2204
rect 11122 2148 11178 2204
rect 11178 2148 11182 2204
rect 11118 2144 11182 2148
rect 11198 2204 11262 2208
rect 11198 2148 11202 2204
rect 11202 2148 11258 2204
rect 11258 2148 11262 2204
rect 11198 2144 11262 2148
rect 11278 2204 11342 2208
rect 11278 2148 11282 2204
rect 11282 2148 11338 2204
rect 11338 2148 11342 2204
rect 11278 2144 11342 2148
rect 11358 2204 11422 2208
rect 11358 2148 11362 2204
rect 11362 2148 11418 2204
rect 11418 2148 11422 2204
rect 11358 2144 11422 2148
rect 17895 2204 17959 2208
rect 17895 2148 17899 2204
rect 17899 2148 17955 2204
rect 17955 2148 17959 2204
rect 17895 2144 17959 2148
rect 17975 2204 18039 2208
rect 17975 2148 17979 2204
rect 17979 2148 18035 2204
rect 18035 2148 18039 2204
rect 17975 2144 18039 2148
rect 18055 2204 18119 2208
rect 18055 2148 18059 2204
rect 18059 2148 18115 2204
rect 18115 2148 18119 2204
rect 18055 2144 18119 2148
rect 18135 2204 18199 2208
rect 18135 2148 18139 2204
rect 18139 2148 18195 2204
rect 18195 2148 18199 2204
rect 18135 2144 18199 2148
<< metal4 >>
rect 4332 21792 4653 22352
rect 4332 21728 4340 21792
rect 4404 21728 4420 21792
rect 4484 21728 4500 21792
rect 4564 21728 4580 21792
rect 4644 21728 4653 21792
rect 4332 20704 4653 21728
rect 4332 20640 4340 20704
rect 4404 20640 4420 20704
rect 4484 20640 4500 20704
rect 4564 20640 4580 20704
rect 4644 20640 4653 20704
rect 4332 19616 4653 20640
rect 4332 19552 4340 19616
rect 4404 19552 4420 19616
rect 4484 19552 4500 19616
rect 4564 19552 4580 19616
rect 4644 19552 4653 19616
rect 4332 19019 4653 19552
rect 4332 18783 4374 19019
rect 4610 18783 4653 19019
rect 4332 18528 4653 18783
rect 4332 18464 4340 18528
rect 4404 18464 4420 18528
rect 4484 18464 4500 18528
rect 4564 18464 4580 18528
rect 4644 18464 4653 18528
rect 4332 17440 4653 18464
rect 4332 17376 4340 17440
rect 4404 17376 4420 17440
rect 4484 17376 4500 17440
rect 4564 17376 4580 17440
rect 4644 17376 4653 17440
rect 4332 16352 4653 17376
rect 4332 16288 4340 16352
rect 4404 16288 4420 16352
rect 4484 16288 4500 16352
rect 4564 16288 4580 16352
rect 4644 16288 4653 16352
rect 4332 15264 4653 16288
rect 4332 15200 4340 15264
rect 4404 15200 4420 15264
rect 4484 15200 4500 15264
rect 4564 15200 4580 15264
rect 4644 15200 4653 15264
rect 4332 14176 4653 15200
rect 4332 14112 4340 14176
rect 4404 14112 4420 14176
rect 4484 14112 4500 14176
rect 4564 14112 4580 14176
rect 4644 14112 4653 14176
rect 4332 13088 4653 14112
rect 4332 13024 4340 13088
rect 4404 13024 4420 13088
rect 4484 13024 4500 13088
rect 4564 13024 4580 13088
rect 4644 13024 4653 13088
rect 4332 12310 4653 13024
rect 4332 12074 4374 12310
rect 4610 12074 4653 12310
rect 4332 12000 4653 12074
rect 4332 11936 4340 12000
rect 4404 11936 4420 12000
rect 4484 11936 4500 12000
rect 4564 11936 4580 12000
rect 4644 11936 4653 12000
rect 4332 10912 4653 11936
rect 4332 10848 4340 10912
rect 4404 10848 4420 10912
rect 4484 10848 4500 10912
rect 4564 10848 4580 10912
rect 4644 10848 4653 10912
rect 4332 9824 4653 10848
rect 4332 9760 4340 9824
rect 4404 9760 4420 9824
rect 4484 9760 4500 9824
rect 4564 9760 4580 9824
rect 4644 9760 4653 9824
rect 4332 8736 4653 9760
rect 4332 8672 4340 8736
rect 4404 8672 4420 8736
rect 4484 8672 4500 8736
rect 4564 8672 4580 8736
rect 4644 8672 4653 8736
rect 4332 7648 4653 8672
rect 4332 7584 4340 7648
rect 4404 7584 4420 7648
rect 4484 7584 4500 7648
rect 4564 7584 4580 7648
rect 4644 7584 4653 7648
rect 4332 6560 4653 7584
rect 4332 6496 4340 6560
rect 4404 6496 4420 6560
rect 4484 6496 4500 6560
rect 4564 6496 4580 6560
rect 4644 6496 4653 6560
rect 4332 5600 4653 6496
rect 4332 5472 4374 5600
rect 4610 5472 4653 5600
rect 4332 5408 4340 5472
rect 4644 5408 4653 5472
rect 4332 5364 4374 5408
rect 4610 5364 4653 5408
rect 4332 4384 4653 5364
rect 4332 4320 4340 4384
rect 4404 4320 4420 4384
rect 4484 4320 4500 4384
rect 4564 4320 4580 4384
rect 4644 4320 4653 4384
rect 4332 3296 4653 4320
rect 4332 3232 4340 3296
rect 4404 3232 4420 3296
rect 4484 3232 4500 3296
rect 4564 3232 4580 3296
rect 4644 3232 4653 3296
rect 4332 2208 4653 3232
rect 4332 2144 4340 2208
rect 4404 2144 4420 2208
rect 4484 2144 4500 2208
rect 4564 2144 4580 2208
rect 4644 2144 4653 2208
rect 4332 2128 4653 2144
rect 7721 22336 8041 22352
rect 7721 22272 7729 22336
rect 7793 22272 7809 22336
rect 7873 22272 7889 22336
rect 7953 22272 7969 22336
rect 8033 22272 8041 22336
rect 7721 21248 8041 22272
rect 7721 21184 7729 21248
rect 7793 21184 7809 21248
rect 7873 21184 7889 21248
rect 7953 21184 7969 21248
rect 8033 21184 8041 21248
rect 7721 20160 8041 21184
rect 7721 20096 7729 20160
rect 7793 20096 7809 20160
rect 7873 20096 7889 20160
rect 7953 20096 7969 20160
rect 8033 20096 8041 20160
rect 7721 19072 8041 20096
rect 7721 19008 7729 19072
rect 7793 19008 7809 19072
rect 7873 19008 7889 19072
rect 7953 19008 7969 19072
rect 8033 19008 8041 19072
rect 7721 17984 8041 19008
rect 7721 17920 7729 17984
rect 7793 17920 7809 17984
rect 7873 17920 7889 17984
rect 7953 17920 7969 17984
rect 8033 17920 8041 17984
rect 7721 16896 8041 17920
rect 7721 16832 7729 16896
rect 7793 16832 7809 16896
rect 7873 16832 7889 16896
rect 7953 16832 7969 16896
rect 8033 16832 8041 16896
rect 7721 15808 8041 16832
rect 7721 15744 7729 15808
rect 7793 15744 7809 15808
rect 7873 15744 7889 15808
rect 7953 15744 7969 15808
rect 8033 15744 8041 15808
rect 7721 15664 8041 15744
rect 7721 15428 7763 15664
rect 7999 15428 8041 15664
rect 7721 14720 8041 15428
rect 7721 14656 7729 14720
rect 7793 14656 7809 14720
rect 7873 14656 7889 14720
rect 7953 14656 7969 14720
rect 8033 14656 8041 14720
rect 7721 13632 8041 14656
rect 7721 13568 7729 13632
rect 7793 13568 7809 13632
rect 7873 13568 7889 13632
rect 7953 13568 7969 13632
rect 8033 13568 8041 13632
rect 7721 12544 8041 13568
rect 7721 12480 7729 12544
rect 7793 12480 7809 12544
rect 7873 12480 7889 12544
rect 7953 12480 7969 12544
rect 8033 12480 8041 12544
rect 7721 11456 8041 12480
rect 7721 11392 7729 11456
rect 7793 11392 7809 11456
rect 7873 11392 7889 11456
rect 7953 11392 7969 11456
rect 8033 11392 8041 11456
rect 7721 10368 8041 11392
rect 7721 10304 7729 10368
rect 7793 10304 7809 10368
rect 7873 10304 7889 10368
rect 7953 10304 7969 10368
rect 8033 10304 8041 10368
rect 7721 9280 8041 10304
rect 7721 9216 7729 9280
rect 7793 9216 7809 9280
rect 7873 9216 7889 9280
rect 7953 9216 7969 9280
rect 8033 9216 8041 9280
rect 7721 8955 8041 9216
rect 7721 8719 7763 8955
rect 7999 8719 8041 8955
rect 7721 8192 8041 8719
rect 7721 8128 7729 8192
rect 7793 8128 7809 8192
rect 7873 8128 7889 8192
rect 7953 8128 7969 8192
rect 8033 8128 8041 8192
rect 7721 7104 8041 8128
rect 7721 7040 7729 7104
rect 7793 7040 7809 7104
rect 7873 7040 7889 7104
rect 7953 7040 7969 7104
rect 8033 7040 8041 7104
rect 7721 6016 8041 7040
rect 7721 5952 7729 6016
rect 7793 5952 7809 6016
rect 7873 5952 7889 6016
rect 7953 5952 7969 6016
rect 8033 5952 8041 6016
rect 7721 4928 8041 5952
rect 7721 4864 7729 4928
rect 7793 4864 7809 4928
rect 7873 4864 7889 4928
rect 7953 4864 7969 4928
rect 8033 4864 8041 4928
rect 7721 3840 8041 4864
rect 7721 3776 7729 3840
rect 7793 3776 7809 3840
rect 7873 3776 7889 3840
rect 7953 3776 7969 3840
rect 8033 3776 8041 3840
rect 7721 2752 8041 3776
rect 7721 2688 7729 2752
rect 7793 2688 7809 2752
rect 7873 2688 7889 2752
rect 7953 2688 7969 2752
rect 8033 2688 8041 2752
rect 7721 2128 8041 2688
rect 11110 21792 11430 22352
rect 11110 21728 11118 21792
rect 11182 21728 11198 21792
rect 11262 21728 11278 21792
rect 11342 21728 11358 21792
rect 11422 21728 11430 21792
rect 11110 20704 11430 21728
rect 11110 20640 11118 20704
rect 11182 20640 11198 20704
rect 11262 20640 11278 20704
rect 11342 20640 11358 20704
rect 11422 20640 11430 20704
rect 11110 19616 11430 20640
rect 11110 19552 11118 19616
rect 11182 19552 11198 19616
rect 11262 19552 11278 19616
rect 11342 19552 11358 19616
rect 11422 19552 11430 19616
rect 11110 19019 11430 19552
rect 11110 18783 11152 19019
rect 11388 18783 11430 19019
rect 11110 18528 11430 18783
rect 11110 18464 11118 18528
rect 11182 18464 11198 18528
rect 11262 18464 11278 18528
rect 11342 18464 11358 18528
rect 11422 18464 11430 18528
rect 11110 17440 11430 18464
rect 11110 17376 11118 17440
rect 11182 17376 11198 17440
rect 11262 17376 11278 17440
rect 11342 17376 11358 17440
rect 11422 17376 11430 17440
rect 11110 16352 11430 17376
rect 11110 16288 11118 16352
rect 11182 16288 11198 16352
rect 11262 16288 11278 16352
rect 11342 16288 11358 16352
rect 11422 16288 11430 16352
rect 11110 15264 11430 16288
rect 11110 15200 11118 15264
rect 11182 15200 11198 15264
rect 11262 15200 11278 15264
rect 11342 15200 11358 15264
rect 11422 15200 11430 15264
rect 11110 14176 11430 15200
rect 11110 14112 11118 14176
rect 11182 14112 11198 14176
rect 11262 14112 11278 14176
rect 11342 14112 11358 14176
rect 11422 14112 11430 14176
rect 11110 13088 11430 14112
rect 11110 13024 11118 13088
rect 11182 13024 11198 13088
rect 11262 13024 11278 13088
rect 11342 13024 11358 13088
rect 11422 13024 11430 13088
rect 11110 12310 11430 13024
rect 11110 12074 11152 12310
rect 11388 12074 11430 12310
rect 11110 12000 11430 12074
rect 11110 11936 11118 12000
rect 11182 11936 11198 12000
rect 11262 11936 11278 12000
rect 11342 11936 11358 12000
rect 11422 11936 11430 12000
rect 11110 10912 11430 11936
rect 11110 10848 11118 10912
rect 11182 10848 11198 10912
rect 11262 10848 11278 10912
rect 11342 10848 11358 10912
rect 11422 10848 11430 10912
rect 11110 9824 11430 10848
rect 11110 9760 11118 9824
rect 11182 9760 11198 9824
rect 11262 9760 11278 9824
rect 11342 9760 11358 9824
rect 11422 9760 11430 9824
rect 11110 8736 11430 9760
rect 11110 8672 11118 8736
rect 11182 8672 11198 8736
rect 11262 8672 11278 8736
rect 11342 8672 11358 8736
rect 11422 8672 11430 8736
rect 11110 7648 11430 8672
rect 11110 7584 11118 7648
rect 11182 7584 11198 7648
rect 11262 7584 11278 7648
rect 11342 7584 11358 7648
rect 11422 7584 11430 7648
rect 11110 6560 11430 7584
rect 11110 6496 11118 6560
rect 11182 6496 11198 6560
rect 11262 6496 11278 6560
rect 11342 6496 11358 6560
rect 11422 6496 11430 6560
rect 11110 5600 11430 6496
rect 11110 5472 11152 5600
rect 11388 5472 11430 5600
rect 11110 5408 11118 5472
rect 11422 5408 11430 5472
rect 11110 5364 11152 5408
rect 11388 5364 11430 5408
rect 11110 4384 11430 5364
rect 11110 4320 11118 4384
rect 11182 4320 11198 4384
rect 11262 4320 11278 4384
rect 11342 4320 11358 4384
rect 11422 4320 11430 4384
rect 11110 3296 11430 4320
rect 11110 3232 11118 3296
rect 11182 3232 11198 3296
rect 11262 3232 11278 3296
rect 11342 3232 11358 3296
rect 11422 3232 11430 3296
rect 11110 2208 11430 3232
rect 11110 2144 11118 2208
rect 11182 2144 11198 2208
rect 11262 2144 11278 2208
rect 11342 2144 11358 2208
rect 11422 2144 11430 2208
rect 11110 2128 11430 2144
rect 14498 22336 14819 22352
rect 14498 22272 14506 22336
rect 14570 22272 14586 22336
rect 14650 22272 14666 22336
rect 14730 22272 14746 22336
rect 14810 22272 14819 22336
rect 14498 21248 14819 22272
rect 14498 21184 14506 21248
rect 14570 21184 14586 21248
rect 14650 21184 14666 21248
rect 14730 21184 14746 21248
rect 14810 21184 14819 21248
rect 14498 20160 14819 21184
rect 14498 20096 14506 20160
rect 14570 20096 14586 20160
rect 14650 20096 14666 20160
rect 14730 20096 14746 20160
rect 14810 20096 14819 20160
rect 14498 19072 14819 20096
rect 14498 19008 14506 19072
rect 14570 19008 14586 19072
rect 14650 19008 14666 19072
rect 14730 19008 14746 19072
rect 14810 19008 14819 19072
rect 14498 17984 14819 19008
rect 14498 17920 14506 17984
rect 14570 17920 14586 17984
rect 14650 17920 14666 17984
rect 14730 17920 14746 17984
rect 14810 17920 14819 17984
rect 14498 16896 14819 17920
rect 14498 16832 14506 16896
rect 14570 16832 14586 16896
rect 14650 16832 14666 16896
rect 14730 16832 14746 16896
rect 14810 16832 14819 16896
rect 14498 15808 14819 16832
rect 14498 15744 14506 15808
rect 14570 15744 14586 15808
rect 14650 15744 14666 15808
rect 14730 15744 14746 15808
rect 14810 15744 14819 15808
rect 14498 15664 14819 15744
rect 14498 15428 14540 15664
rect 14776 15428 14819 15664
rect 14498 14720 14819 15428
rect 14498 14656 14506 14720
rect 14570 14656 14586 14720
rect 14650 14656 14666 14720
rect 14730 14656 14746 14720
rect 14810 14656 14819 14720
rect 14498 13632 14819 14656
rect 14498 13568 14506 13632
rect 14570 13568 14586 13632
rect 14650 13568 14666 13632
rect 14730 13568 14746 13632
rect 14810 13568 14819 13632
rect 14498 12544 14819 13568
rect 14498 12480 14506 12544
rect 14570 12480 14586 12544
rect 14650 12480 14666 12544
rect 14730 12480 14746 12544
rect 14810 12480 14819 12544
rect 14498 11456 14819 12480
rect 14498 11392 14506 11456
rect 14570 11392 14586 11456
rect 14650 11392 14666 11456
rect 14730 11392 14746 11456
rect 14810 11392 14819 11456
rect 14498 10368 14819 11392
rect 14498 10304 14506 10368
rect 14570 10304 14586 10368
rect 14650 10304 14666 10368
rect 14730 10304 14746 10368
rect 14810 10304 14819 10368
rect 14498 9280 14819 10304
rect 14498 9216 14506 9280
rect 14570 9216 14586 9280
rect 14650 9216 14666 9280
rect 14730 9216 14746 9280
rect 14810 9216 14819 9280
rect 14498 8955 14819 9216
rect 14498 8719 14540 8955
rect 14776 8719 14819 8955
rect 14498 8192 14819 8719
rect 14498 8128 14506 8192
rect 14570 8128 14586 8192
rect 14650 8128 14666 8192
rect 14730 8128 14746 8192
rect 14810 8128 14819 8192
rect 14498 7104 14819 8128
rect 14498 7040 14506 7104
rect 14570 7040 14586 7104
rect 14650 7040 14666 7104
rect 14730 7040 14746 7104
rect 14810 7040 14819 7104
rect 14498 6016 14819 7040
rect 14498 5952 14506 6016
rect 14570 5952 14586 6016
rect 14650 5952 14666 6016
rect 14730 5952 14746 6016
rect 14810 5952 14819 6016
rect 14498 4928 14819 5952
rect 14498 4864 14506 4928
rect 14570 4864 14586 4928
rect 14650 4864 14666 4928
rect 14730 4864 14746 4928
rect 14810 4864 14819 4928
rect 14498 3840 14819 4864
rect 14498 3776 14506 3840
rect 14570 3776 14586 3840
rect 14650 3776 14666 3840
rect 14730 3776 14746 3840
rect 14810 3776 14819 3840
rect 14498 2752 14819 3776
rect 14498 2688 14506 2752
rect 14570 2688 14586 2752
rect 14650 2688 14666 2752
rect 14730 2688 14746 2752
rect 14810 2688 14819 2752
rect 14498 2128 14819 2688
rect 17887 21792 18207 22352
rect 17887 21728 17895 21792
rect 17959 21728 17975 21792
rect 18039 21728 18055 21792
rect 18119 21728 18135 21792
rect 18199 21728 18207 21792
rect 17887 20704 18207 21728
rect 17887 20640 17895 20704
rect 17959 20640 17975 20704
rect 18039 20640 18055 20704
rect 18119 20640 18135 20704
rect 18199 20640 18207 20704
rect 17887 19616 18207 20640
rect 17887 19552 17895 19616
rect 17959 19552 17975 19616
rect 18039 19552 18055 19616
rect 18119 19552 18135 19616
rect 18199 19552 18207 19616
rect 17887 19019 18207 19552
rect 17887 18783 17929 19019
rect 18165 18783 18207 19019
rect 17887 18528 18207 18783
rect 17887 18464 17895 18528
rect 17959 18464 17975 18528
rect 18039 18464 18055 18528
rect 18119 18464 18135 18528
rect 18199 18464 18207 18528
rect 17887 17440 18207 18464
rect 17887 17376 17895 17440
rect 17959 17376 17975 17440
rect 18039 17376 18055 17440
rect 18119 17376 18135 17440
rect 18199 17376 18207 17440
rect 17887 16352 18207 17376
rect 17887 16288 17895 16352
rect 17959 16288 17975 16352
rect 18039 16288 18055 16352
rect 18119 16288 18135 16352
rect 18199 16288 18207 16352
rect 17887 15264 18207 16288
rect 17887 15200 17895 15264
rect 17959 15200 17975 15264
rect 18039 15200 18055 15264
rect 18119 15200 18135 15264
rect 18199 15200 18207 15264
rect 17887 14176 18207 15200
rect 17887 14112 17895 14176
rect 17959 14112 17975 14176
rect 18039 14112 18055 14176
rect 18119 14112 18135 14176
rect 18199 14112 18207 14176
rect 17887 13088 18207 14112
rect 17887 13024 17895 13088
rect 17959 13024 17975 13088
rect 18039 13024 18055 13088
rect 18119 13024 18135 13088
rect 18199 13024 18207 13088
rect 17887 12310 18207 13024
rect 17887 12074 17929 12310
rect 18165 12074 18207 12310
rect 17887 12000 18207 12074
rect 17887 11936 17895 12000
rect 17959 11936 17975 12000
rect 18039 11936 18055 12000
rect 18119 11936 18135 12000
rect 18199 11936 18207 12000
rect 17887 10912 18207 11936
rect 17887 10848 17895 10912
rect 17959 10848 17975 10912
rect 18039 10848 18055 10912
rect 18119 10848 18135 10912
rect 18199 10848 18207 10912
rect 17887 9824 18207 10848
rect 17887 9760 17895 9824
rect 17959 9760 17975 9824
rect 18039 9760 18055 9824
rect 18119 9760 18135 9824
rect 18199 9760 18207 9824
rect 17887 8736 18207 9760
rect 17887 8672 17895 8736
rect 17959 8672 17975 8736
rect 18039 8672 18055 8736
rect 18119 8672 18135 8736
rect 18199 8672 18207 8736
rect 17887 7648 18207 8672
rect 17887 7584 17895 7648
rect 17959 7584 17975 7648
rect 18039 7584 18055 7648
rect 18119 7584 18135 7648
rect 18199 7584 18207 7648
rect 17887 6560 18207 7584
rect 17887 6496 17895 6560
rect 17959 6496 17975 6560
rect 18039 6496 18055 6560
rect 18119 6496 18135 6560
rect 18199 6496 18207 6560
rect 17887 5600 18207 6496
rect 17887 5472 17929 5600
rect 18165 5472 18207 5600
rect 17887 5408 17895 5472
rect 18199 5408 18207 5472
rect 17887 5364 17929 5408
rect 18165 5364 18207 5408
rect 17887 4384 18207 5364
rect 17887 4320 17895 4384
rect 17959 4320 17975 4384
rect 18039 4320 18055 4384
rect 18119 4320 18135 4384
rect 18199 4320 18207 4384
rect 17887 3296 18207 4320
rect 17887 3232 17895 3296
rect 17959 3232 17975 3296
rect 18039 3232 18055 3296
rect 18119 3232 18135 3296
rect 18199 3232 18207 3296
rect 17887 2208 18207 3232
rect 17887 2144 17895 2208
rect 17959 2144 17975 2208
rect 18039 2144 18055 2208
rect 18119 2144 18135 2208
rect 18199 2144 18207 2208
rect 17887 2128 18207 2144
<< via4 >>
rect 4374 18783 4610 19019
rect 4374 12074 4610 12310
rect 4374 5472 4610 5600
rect 4374 5408 4404 5472
rect 4404 5408 4420 5472
rect 4420 5408 4484 5472
rect 4484 5408 4500 5472
rect 4500 5408 4564 5472
rect 4564 5408 4580 5472
rect 4580 5408 4610 5472
rect 4374 5364 4610 5408
rect 7763 15428 7999 15664
rect 7763 8719 7999 8955
rect 11152 18783 11388 19019
rect 11152 12074 11388 12310
rect 11152 5472 11388 5600
rect 11152 5408 11182 5472
rect 11182 5408 11198 5472
rect 11198 5408 11262 5472
rect 11262 5408 11278 5472
rect 11278 5408 11342 5472
rect 11342 5408 11358 5472
rect 11358 5408 11388 5472
rect 11152 5364 11388 5408
rect 14540 15428 14776 15664
rect 14540 8719 14776 8955
rect 17929 18783 18165 19019
rect 17929 12074 18165 12310
rect 17929 5472 18165 5600
rect 17929 5408 17959 5472
rect 17959 5408 17975 5472
rect 17975 5408 18039 5472
rect 18039 5408 18055 5472
rect 18055 5408 18119 5472
rect 18119 5408 18135 5472
rect 18135 5408 18165 5472
rect 17929 5364 18165 5408
<< metal5 >>
rect 1104 19019 21436 19061
rect 1104 18783 4374 19019
rect 4610 18783 11152 19019
rect 11388 18783 17929 19019
rect 18165 18783 21436 19019
rect 1104 18741 21436 18783
rect 1104 15664 21436 15707
rect 1104 15428 7763 15664
rect 7999 15428 14540 15664
rect 14776 15428 21436 15664
rect 1104 15386 21436 15428
rect 1104 12310 21436 12352
rect 1104 12074 4374 12310
rect 4610 12074 11152 12310
rect 11388 12074 17929 12310
rect 18165 12074 21436 12310
rect 1104 12032 21436 12074
rect 1104 8955 21436 8997
rect 1104 8719 7763 8955
rect 7999 8719 14540 8955
rect 14776 8719 21436 8955
rect 1104 8677 21436 8719
rect 1104 5600 21436 5643
rect 1104 5364 4374 5600
rect 4610 5364 11152 5600
rect 11388 5364 17929 5600
rect 18165 5364 21436 5600
rect 1104 5322 21436 5364
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1617727139
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1617727139
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1617727139
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1617727139
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1617727139
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1617727139
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 1617727139
transform 1 0 4324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1617727139
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1617727139
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1617727139
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1617727139
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _131_
timestamp 1617727139
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1617727139
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1617727139
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_45
timestamp 1617727139
transform 1 0 5244 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1617727139
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1617727139
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1617727139
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1617727139
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1617727139
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82
timestamp 1617727139
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_70
timestamp 1617727139
transform 1 0 7544 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _111_
timestamp 1617727139
transform 1 0 6900 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1617727139
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1617727139
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94
timestamp 1617727139
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1617727139
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1617727139
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _112_
timestamp 1617727139
transform 1 0 10488 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1617727139
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1617727139
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1617727139
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1617727139
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114
timestamp 1617727139
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1617727139
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1617727139
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1617727139
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1617727139
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1617727139
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1617727139
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1617727139
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1617727139
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1617727139
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1617727139
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1617727139
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1617727139
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1617727139
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1617727139
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1617727139
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1617727139
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1617727139
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_196
timestamp 1617727139
transform 1 0 19136 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1617727139
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1617727139
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_210
timestamp 1617727139
transform 1 0 20424 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1617727139
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1617727139
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1617727139
transform -1 0 21436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1617727139
transform -1 0 21436 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1617727139
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1617727139
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1617727139
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1617727139
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1617727139
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1617727139
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1617727139
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1617727139
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1617727139
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1617727139
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_101
timestamp 1617727139
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1617727139
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1617727139
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1617727139
transform 1 0 10672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_119
timestamp 1617727139
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_107
timestamp 1617727139
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_143
timestamp 1617727139
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_131
timestamp 1617727139
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1617727139
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1617727139
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1617727139
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1617727139
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1617727139
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1617727139
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1617727139
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_215
timestamp 1617727139
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1617727139
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1617727139
transform -1 0 21436 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1617727139
transform 1 0 2484 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1617727139
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1617727139
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_36
timestamp 1617727139
transform 1 0 4416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_21
timestamp 1617727139
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _099_
timestamp 1617727139
transform 1 0 3128 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1617727139
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1617727139
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_48
timestamp 1617727139
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1617727139
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1617727139
transform 1 0 8556 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1617727139
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _147_
timestamp 1617727139
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1617727139
transform 1 0 9660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1617727139
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1617727139
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1617727139
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1617727139
transform 1 0 10764 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1617727139
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _149_
timestamp 1617727139
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_145
timestamp 1617727139
transform 1 0 14444 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_133
timestamp 1617727139
transform 1 0 13340 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_157
timestamp 1617727139
transform 1 0 15548 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1617727139
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1617727139
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1617727139
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1617727139
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_208
timestamp 1617727139
transform 1 0 20240 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1617727139
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_216
timestamp 1617727139
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1617727139
transform -1 0 21436 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_18
timestamp 1617727139
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_6
timestamp 1617727139
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1617727139
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1617727139
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1617727139
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1617727139
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1617727139
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1617727139
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _106_
timestamp 1617727139
transform 1 0 6256 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1617727139
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_69
timestamp 1617727139
transform 1 0 7452 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1617727139
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1617727139
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1617727139
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1617727139
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1617727139
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1617727139
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1617727139
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_160
timestamp 1617727139
transform 1 0 15824 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1617727139
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1617727139
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _154_
timestamp 1617727139
transform 1 0 15916 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1617727139
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_204
timestamp 1617727139
transform 1 0 19872 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_192
timestamp 1617727139
transform 1 0 18768 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp 1617727139
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1617727139
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1617727139
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1617727139
transform -1 0 21436 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1617727139
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1617727139
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1617727139
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1617727139
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1617727139
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1617727139
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1617727139
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1617727139
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1617727139
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1617727139
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1617727139
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1617727139
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1617727139
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1617727139
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1617727139
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1617727139
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1617727139
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1617727139
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1617727139
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1617727139
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1617727139
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_208
timestamp 1617727139
transform 1 0 20240 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1617727139
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1617727139
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1617727139
transform -1 0 21436 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1617727139
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1617727139
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11
timestamp 1617727139
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1617727139
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1617727139
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1617727139
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _130_
timestamp 1617727139
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _109_
timestamp 1617727139
transform 1 0 2300 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_37
timestamp 1617727139
transform 1 0 4508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_25
timestamp 1617727139
transform 1 0 3404 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1617727139
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1617727139
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1617727139
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1617727139
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_49
timestamp 1617727139
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1617727139
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1617727139
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1617727139
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1617727139
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1617727139
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1617727139
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1617727139
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1617727139
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1617727139
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1617727139
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1617727139
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1617727139
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1617727139
transform 1 0 11684 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 1617727139
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1617727139
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _141_
timestamp 1617727139
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1617727139
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1617727139
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1617727139
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1617727139
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1617727139
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1617727139
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1617727139
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1617727139
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1617727139
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1617727139
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1617727139
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1617727139
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1617727139
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_208
timestamp 1617727139
transform 1 0 20240 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1617727139
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1617727139
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1617727139
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1617727139
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp 1617727139
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1617727139
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1617727139
transform -1 0 21436 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1617727139
transform -1 0 21436 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_19
timestamp 1617727139
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1617727139
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1617727139
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1617727139
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _082_
timestamp 1617727139
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1617727139
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1617727139
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1617727139
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1617727139
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1617727139
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _151_
timestamp 1617727139
transform 1 0 6992 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1617727139
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_93
timestamp 1617727139
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1617727139
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1617727139
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1617727139
transform 1 0 10212 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_114
timestamp 1617727139
transform 1 0 11592 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_138
timestamp 1617727139
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_126
timestamp 1617727139
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1617727139
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1617727139
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1617727139
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _083_
timestamp 1617727139
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_187
timestamp 1617727139
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1617727139
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_206
timestamp 1617727139
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _115_
timestamp 1617727139
transform 1 0 19412 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1617727139
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1617727139
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1617727139
transform -1 0 21436 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1617727139
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1617727139
transform 1 0 1748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1617727139
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1617727139
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1617727139
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_4  _140_
timestamp 1617727139
transform 1 0 3036 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1617727139
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1617727139
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1617727139
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1617727139
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1617727139
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1617727139
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_86
timestamp 1617727139
transform 1 0 9016 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _097_
timestamp 1617727139
transform 1 0 9568 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1617727139
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1617727139
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_111
timestamp 1617727139
transform 1 0 11316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1617727139
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1617727139
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_160
timestamp 1617727139
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_147
timestamp 1617727139
transform 1 0 14628 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _089_
timestamp 1617727139
transform 1 0 15180 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1617727139
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1617727139
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1617727139
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1617727139
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_208
timestamp 1617727139
transform 1 0 20240 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1617727139
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1617727139
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1617727139
transform -1 0 21436 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_17
timestamp 1617727139
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1617727139
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1617727139
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1617727139
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1617727139
transform 1 0 2392 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1617727139
transform 1 0 4692 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1617727139
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1617727139
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _114_
timestamp 1617727139
transform 1 0 4048 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_51
timestamp 1617727139
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_75
timestamp 1617727139
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_63
timestamp 1617727139
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1617727139
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1617727139
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1617727139
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1617727139
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1617727139
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1617727139
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1617727139
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1617727139
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1617727139
transform 1 0 16376 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1617727139
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1617727139
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1617727139
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1617727139
transform 1 0 16744 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _113_
timestamp 1617727139
transform 1 0 16836 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1617727139
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_192
timestamp 1617727139
transform 1 0 18768 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1617727139
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1617727139
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1617727139
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1617727139
transform -1 0 21436 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1617727139
transform 1 0 2484 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1617727139
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1617727139
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1617727139
transform 1 0 4876 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1617727139
transform 1 0 3772 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_23
timestamp 1617727139
transform 1 0 3220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1617727139
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1617727139
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1617727139
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1617727139
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_83
timestamp 1617727139
transform 1 0 8740 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _160_
timestamp 1617727139
transform 1 0 6992 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_95
timestamp 1617727139
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1617727139
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1617727139
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_107
timestamp 1617727139
transform 1 0 10948 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1617727139
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1617727139
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_162
timestamp 1617727139
transform 1 0 16008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_147
timestamp 1617727139
transform 1 0 14628 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _136_
timestamp 1617727139
transform 1 0 15180 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1617727139
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1617727139
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1617727139
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1617727139
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_208
timestamp 1617727139
transform 1 0 20240 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1617727139
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1617727139
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1617727139
transform -1 0 21436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1617727139
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _157_
timestamp 1617727139
transform 1 0 1380 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1617727139
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1617727139
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1617727139
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1617727139
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1617727139
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1617727139
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1617727139
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1617727139
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_101
timestamp 1617727139
transform 1 0 10396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1617727139
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1617727139
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _095_
timestamp 1617727139
transform 1 0 9752 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_124
timestamp 1617727139
transform 1 0 12512 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_112
timestamp 1617727139
transform 1 0 11408 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1617727139
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1617727139
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _134_
timestamp 1617727139
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1617727139
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1617727139
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1617727139
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1617727139
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1617727139
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1617727139
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_215
timestamp 1617727139
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1617727139
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1617727139
transform -1 0 21436 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1617727139
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1617727139
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1617727139
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1617727139
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1617727139
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1617727139
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _119_
timestamp 1617727139
transform 1 0 1656 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1617727139
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1617727139
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1617727139
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1617727139
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1617727139
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1617727139
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1617727139
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1617727139
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1617727139
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1617727139
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1617727139
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1617727139
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1617727139
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1617727139
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_74
timestamp 1617727139
transform 1 0 7912 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1617727139
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1617727139
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1617727139
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1617727139
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1617727139
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1617727139
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _123_
timestamp 1617727139
transform 1 0 10120 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1617727139
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1617727139
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1617727139
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1617727139
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1617727139
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1617727139
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1617727139
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1617727139
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1617727139
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1617727139
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1617727139
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1617727139
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1617727139
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1617727139
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1617727139
transform 1 0 17388 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1617727139
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1617727139
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1617727139
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _138_
timestamp 1617727139
transform 1 0 16560 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1617727139
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_189
timestamp 1617727139
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_204
timestamp 1617727139
transform 1 0 19872 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_196
timestamp 1617727139
transform 1 0 19136 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _142_
timestamp 1617727139
transform 1 0 18768 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1617727139
transform 1 0 19964 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_215
timestamp 1617727139
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1617727139
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_217
timestamp 1617727139
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_209
timestamp 1617727139
transform 1 0 20332 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1617727139
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1617727139
transform -1 0 21436 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1617727139
transform -1 0 21436 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1617727139
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1617727139
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1617727139
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1617727139
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1617727139
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1617727139
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1617727139
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1617727139
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1617727139
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1617727139
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_72
timestamp 1617727139
transform 1 0 7728 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _146_
timestamp 1617727139
transform 1 0 7084 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _137_
timestamp 1617727139
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_103
timestamp 1617727139
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_91
timestamp 1617727139
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1617727139
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1617727139
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1617727139
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1617727139
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1617727139
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _155_
timestamp 1617727139
transform 1 0 12880 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1617727139
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1617727139
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _102_
timestamp 1617727139
transform 1 0 16100 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1617727139
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1617727139
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_170
timestamp 1617727139
transform 1 0 16744 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1617727139
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_200
timestamp 1617727139
transform 1 0 19504 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1617727139
transform 1 0 19136 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _117_
timestamp 1617727139
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_210
timestamp 1617727139
transform 1 0 20424 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1617727139
transform -1 0 21436 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1617727139
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1617727139
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1617727139
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1617727139
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1617727139
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1617727139
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _116_
timestamp 1617727139
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1617727139
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1617727139
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _101_
timestamp 1617727139
transform 1 0 6808 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_16_75
timestamp 1617727139
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1617727139
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1617727139
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1617727139
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _159_
timestamp 1617727139
transform 1 0 9660 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_124
timestamp 1617727139
transform 1 0 12512 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_112
timestamp 1617727139
transform 1 0 11408 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_136
timestamp 1617727139
transform 1 0 13616 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1617727139
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1617727139
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1617727139
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1617727139
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1617727139
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1617727139
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1617727139
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1617727139
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 1617727139
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1617727139
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1617727139
transform -1 0 21436 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1617727139
transform 1 0 2484 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1617727139
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1617727139
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1617727139
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_23
timestamp 1617727139
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _100_
timestamp 1617727139
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1617727139
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1617727139
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_47
timestamp 1617727139
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1617727139
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1617727139
transform 1 0 7912 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1617727139
transform 1 0 8648 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_17_102
timestamp 1617727139
transform 1 0 10488 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_114
timestamp 1617727139
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1617727139
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _133_
timestamp 1617727139
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1617727139
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_132
timestamp 1617727139
transform 1 0 13248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_160
timestamp 1617727139
transform 1 0 15824 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1617727139
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _078_
timestamp 1617727139
transform 1 0 15916 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1617727139
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1617727139
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_168
timestamp 1617727139
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1617727139
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_208
timestamp 1617727139
transform 1 0 20240 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1617727139
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1617727139
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1617727139
transform -1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1617727139
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1617727139
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1617727139
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1617727139
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1617727139
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1617727139
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1617727139
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1617727139
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1617727139
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1617727139
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_101
timestamp 1617727139
transform 1 0 10396 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_93
timestamp 1617727139
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1617727139
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _153_
timestamp 1617727139
transform 1 0 10672 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1617727139
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_135
timestamp 1617727139
transform 1 0 13524 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1617727139
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1617727139
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1617727139
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1617727139
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1617727139
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1617727139
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1617727139
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_215
timestamp 1617727139
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1617727139
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1617727139
transform -1 0 21436 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1617727139
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1617727139
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1617727139
transform 1 0 2484 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1617727139
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1617727139
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1617727139
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1617727139
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1617727139
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1617727139
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _150_
timestamp 1617727139
transform 1 0 3220 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1617727139
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1617727139
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1617727139
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1617727139
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_54
timestamp 1617727139
transform 1 0 6072 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1617727139
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1617727139
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1617727139
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1617727139
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1617727139
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1617727139
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1617727139
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1617727139
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1617727139
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1617727139
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1617727139
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1617727139
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1617727139
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1617727139
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1617727139
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1617727139
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1617727139
transform 1 0 14076 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_135
timestamp 1617727139
transform 1 0 13524 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _098_
timestamp 1617727139
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1617727139
transform 1 0 16376 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1617727139
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_163
timestamp 1617727139
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1617727139
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1617727139
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1617727139
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1617727139
transform 1 0 16744 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1617727139
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1617727139
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1617727139
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _085_
timestamp 1617727139
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_204
timestamp 1617727139
transform 1 0 19872 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_192
timestamp 1617727139
transform 1 0 18768 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_200
timestamp 1617727139
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1617727139
transform 1 0 19136 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _126_
timestamp 1617727139
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1617727139
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1617727139
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_210
timestamp 1617727139
transform 1 0 20424 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1617727139
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1617727139
transform -1 0 21436 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1617727139
transform -1 0 21436 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1617727139
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1617727139
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1617727139
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1617727139
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1617727139
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1617727139
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1617727139
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1617727139
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1617727139
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1617727139
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1617727139
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1617727139
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1617727139
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1617727139
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1617727139
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1617727139
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1617727139
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1617727139
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1617727139
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1617727139
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1617727139
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_208
timestamp 1617727139
transform 1 0 20240 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1617727139
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_216
timestamp 1617727139
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1617727139
transform -1 0 21436 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1617727139
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1617727139
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1617727139
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1617727139
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1617727139
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _152_
timestamp 1617727139
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_51
timestamp 1617727139
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_83
timestamp 1617727139
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_79
timestamp 1617727139
transform 1 0 8372 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1617727139
transform 1 0 8004 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1617727139
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1617727139
transform 1 0 8464 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1617727139
transform 1 0 10028 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1617727139
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1617727139
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1617727139
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1617727139
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1617727139
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1617727139
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_133
timestamp 1617727139
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1617727139
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1617727139
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1617727139
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _103_
timestamp 1617727139
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1617727139
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1617727139
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1617727139
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1617727139
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1617727139
transform -1 0 21436 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1617727139
transform 1 0 2484 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1617727139
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1617727139
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1617727139
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _161_
timestamp 1617727139
transform 1 0 3496 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1617727139
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1617727139
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_45
timestamp 1617727139
transform 1 0 5244 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1617727139
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1617727139
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1617727139
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1617727139
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1617727139
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1617727139
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1617727139
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_138
timestamp 1617727139
transform 1 0 13800 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _121_
timestamp 1617727139
transform 1 0 12696 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1617727139
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1617727139
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _139_
timestamp 1617727139
transform 1 0 15088 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1617727139
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1617727139
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1617727139
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_208
timestamp 1617727139
transform 1 0 20240 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1617727139
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_216
timestamp 1617727139
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1617727139
transform -1 0 21436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1617727139
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1617727139
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1617727139
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_32
timestamp 1617727139
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1617727139
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1617727139
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1617727139
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_55
timestamp 1617727139
transform 1 0 6164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_43
timestamp 1617727139
transform 1 0 5060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_79
timestamp 1617727139
transform 1 0 8372 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_67
timestamp 1617727139
transform 1 0 7268 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1617727139
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1617727139
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1617727139
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1617727139
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1617727139
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1617727139
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1617727139
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_157
timestamp 1617727139
transform 1 0 15548 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1617727139
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1617727139
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_181
timestamp 1617727139
transform 1 0 17756 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_169
timestamp 1617727139
transform 1 0 16652 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1617727139
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_193
timestamp 1617727139
transform 1 0 18860 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_215
timestamp 1617727139
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1617727139
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1617727139
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1617727139
transform -1 0 21436 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1617727139
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1617727139
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1617727139
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1617727139
transform 1 0 2852 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_34
timestamp 1617727139
transform 1 0 4232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_22
timestamp 1617727139
transform 1 0 3128 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1617727139
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_46
timestamp 1617727139
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1617727139
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _105_
timestamp 1617727139
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1617727139
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1617727139
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1617727139
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1617727139
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1617727139
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1617727139
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_139
timestamp 1617727139
transform 1 0 13892 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1617727139
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _120_
timestamp 1617727139
transform 1 0 13984 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1617727139
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1617727139
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1617727139
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1617727139
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1617727139
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_208
timestamp 1617727139
transform 1 0 20240 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1617727139
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 1617727139
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1617727139
transform -1 0 21436 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1617727139
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1617727139
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1617727139
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1617727139
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1617727139
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1617727139
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1617727139
transform 1 0 3588 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1617727139
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1617727139
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1617727139
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _087_
timestamp 1617727139
transform 1 0 3864 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1617727139
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_54
timestamp 1617727139
transform 1 0 6072 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1617727139
transform 1 0 4968 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1617727139
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1617727139
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1617727139
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1617727139
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_78
timestamp 1617727139
transform 1 0 8280 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_66
timestamp 1617727139
transform 1 0 7176 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1617727139
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1617727139
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1617727139
transform 1 0 10488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1617727139
transform 1 0 9384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1617727139
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1617727139
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1617727139
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1617727139
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1617727139
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1617727139
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1617727139
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1617727139
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1617727139
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_132
timestamp 1617727139
transform 1 0 13248 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1617727139
transform 1 0 12972 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1617727139
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1617727139
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_162
timestamp 1617727139
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1617727139
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1617727139
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1617727139
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _124_
timestamp 1617727139
transform 1 0 16100 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1617727139
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1617727139
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1617727139
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1617727139
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1617727139
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1617727139
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1617727139
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1617727139
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1617727139
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1617727139
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1617727139
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1617727139
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1617727139
transform -1 0 21436 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1617727139
transform -1 0 21436 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_12
timestamp 1617727139
transform 1 0 2208 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1617727139
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _143_
timestamp 1617727139
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1617727139
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1617727139
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_24
timestamp 1617727139
transform 1 0 3312 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1617727139
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1617727139
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1617727139
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1617727139
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1617727139
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1617727139
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1617727139
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1617727139
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1617727139
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1617727139
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1617727139
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1617727139
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _145_
timestamp 1617727139
transform 1 0 15272 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1617727139
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1617727139
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1617727139
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_192
timestamp 1617727139
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_215
timestamp 1617727139
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1617727139
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1617727139
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1617727139
transform -1 0 21436 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1617727139
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1617727139
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1617727139
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1617727139
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1617727139
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1617727139
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1617727139
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1617727139
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _128_
timestamp 1617727139
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_83
timestamp 1617727139
transform 1 0 8740 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_71
timestamp 1617727139
transform 1 0 7636 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_95
timestamp 1617727139
transform 1 0 9844 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1617727139
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1617727139
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_107
timestamp 1617727139
transform 1 0 10948 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1617727139
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1617727139
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1617727139
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1617727139
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1617727139
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1617727139
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1617727139
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_204
timestamp 1617727139
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_196
timestamp 1617727139
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1617727139
transform 1 0 20056 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_210
timestamp 1617727139
transform 1 0 20424 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1617727139
transform -1 0 21436 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1617727139
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1617727139
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1617727139
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1617727139
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1617727139
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1617727139
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1617727139
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1617727139
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1617727139
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1617727139
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1617727139
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1617727139
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1617727139
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1617727139
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1617727139
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1617727139
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_154
timestamp 1617727139
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1617727139
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _158_
timestamp 1617727139
transform 1 0 15824 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_30_179
timestamp 1617727139
transform 1 0 17572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_203
timestamp 1617727139
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_191
timestamp 1617727139
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_215
timestamp 1617727139
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1617727139
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1617727139
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1617727139
transform -1 0 21436 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_12
timestamp 1617727139
transform 1 0 2208 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1617727139
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1617727139
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1617727139
transform 1 0 1932 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_36
timestamp 1617727139
transform 1 0 4416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_24
timestamp 1617727139
transform 1 0 3312 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_62
timestamp 1617727139
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1617727139
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_48
timestamp 1617727139
transform 1 0 5520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1617727139
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_68
timestamp 1617727139
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _162_
timestamp 1617727139
transform 1 0 7452 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_100
timestamp 1617727139
transform 1 0 10304 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_88
timestamp 1617727139
transform 1 0 9200 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1617727139
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1617727139
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_112
timestamp 1617727139
transform 1 0 11408 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1617727139
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1617727139
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _156_
timestamp 1617727139
transform 1 0 13340 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_164
timestamp 1617727139
transform 1 0 16192 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_152
timestamp 1617727139
transform 1 0 15088 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1617727139
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1617727139
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1617727139
transform 1 0 17296 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1617727139
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_208
timestamp 1617727139
transform 1 0 20240 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1617727139
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1617727139
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1617727139
transform -1 0 21436 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1617727139
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1617727139
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1617727139
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _122_
timestamp 1617727139
transform 1 0 1840 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1617727139
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1617727139
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_22
timestamp 1617727139
transform 1 0 3128 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1617727139
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1617727139
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1617727139
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1617727139
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1617727139
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1617727139
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1617727139
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1617727139
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1617727139
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1617727139
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1617727139
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1617727139
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1617727139
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _093_
timestamp 1617727139
transform 1 0 16376 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_185
timestamp 1617727139
transform 1 0 18124 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_173
timestamp 1617727139
transform 1 0 17020 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1617727139
transform 1 0 19228 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1617727139
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1617727139
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1617727139
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1617727139
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1617727139
transform -1 0 21436 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1617727139
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1617727139
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1617727139
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1617727139
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1617727139
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1617727139
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1617727139
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1617727139
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1617727139
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1617727139
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1617727139
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1617727139
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1617727139
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1617727139
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1617727139
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1617727139
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1617727139
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1617727139
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1617727139
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1617727139
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1617727139
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1617727139
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1617727139
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1617727139
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_117
timestamp 1617727139
transform 1 0 11868 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1617727139
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1617727139
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1617727139
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1617727139
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _107_
timestamp 1617727139
transform 1 0 12420 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_144
timestamp 1617727139
transform 1 0 14352 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_132
timestamp 1617727139
transform 1 0 13248 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_142
timestamp 1617727139
transform 1 0 14168 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1617727139
transform 1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1617727139
transform 1 0 13892 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1617727139
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1617727139
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1617727139
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_166
timestamp 1617727139
transform 1 0 16376 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1617727139
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1617727139
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1617727139
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1617727139
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1617727139
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_174
timestamp 1617727139
transform 1 0 17112 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_170
timestamp 1617727139
transform 1 0 16744 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1617727139
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1617727139
transform 1 0 16836 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1617727139
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1617727139
transform 1 0 18584 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_204
timestamp 1617727139
transform 1 0 19872 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_196
timestamp 1617727139
transform 1 0 19136 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _132_
timestamp 1617727139
transform 1 0 18676 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1617727139
transform 1 0 20148 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_215
timestamp 1617727139
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1617727139
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_210
timestamp 1617727139
transform 1 0 20424 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1617727139
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1617727139
transform -1 0 21436 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1617727139
transform -1 0 21436 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1617727139
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1617727139
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1617727139
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1617727139
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1617727139
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1617727139
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1617727139
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1617727139
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1617727139
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1617727139
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_95
timestamp 1617727139
transform 1 0 9844 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_86
timestamp 1617727139
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _081_
timestamp 1617727139
transform 1 0 9200 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1617727139
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1617727139
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_107
timestamp 1617727139
transform 1 0 10948 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1617727139
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1617727139
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1617727139
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1617727139
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_184
timestamp 1617727139
transform 1 0 18032 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1617727139
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1617727139
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _084_
timestamp 1617727139
transform 1 0 18124 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_194
timestamp 1617727139
transform 1 0 18952 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _118_
timestamp 1617727139
transform 1 0 19688 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_35_217
timestamp 1617727139
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_209
timestamp 1617727139
transform 1 0 20332 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1617727139
transform -1 0 21436 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1617727139
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1617727139
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1617727139
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1617727139
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1617727139
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1617727139
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1617727139
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1617727139
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1617727139
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_75
timestamp 1617727139
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1617727139
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_94
timestamp 1617727139
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_87
timestamp 1617727139
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1617727139
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_125
timestamp 1617727139
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_118
timestamp 1617727139
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_106
timestamp 1617727139
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1617727139
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_137
timestamp 1617727139
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1617727139
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_149
timestamp 1617727139
transform 1 0 14812 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1617727139
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1617727139
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1617727139
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1617727139
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _148_
timestamp 1617727139
transform 1 0 18308 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1617727139
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_194
timestamp 1617727139
transform 1 0 18952 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_214
timestamp 1617727139
transform 1 0 20792 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1617727139
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1617727139
transform -1 0 21436 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal2 s 12898 0 12954 800 4 change[0]
port 1 nsew
rlabel metal2 s 21914 23933 21970 24733 4 change[1]
port 2 nsew
rlabel metal2 s 6642 0 6698 800 4 choice[0]
port 3 nsew
rlabel metal2 s 570 0 626 800 4 choice[1]
port 4 nsew
rlabel metal3 s 21789 14696 22589 14816 4 choice[2]
port 5 nsew
rlabel metal2 s 3330 23933 3386 24733 4 clk
port 6 nsew
rlabel metal3 s 0 9800 800 9920 4 coin[0]
port 7 nsew
rlabel metal2 s 19154 0 19210 800 4 coin[1]
port 8 nsew
rlabel metal3 s 21789 5448 22589 5568 4 out[0]
port 9 nsew
rlabel metal3 s 0 19048 800 19168 4 out[1]
port 10 nsew
rlabel metal2 s 15842 23933 15898 24733 4 out[2]
port 11 nsew
rlabel metal2 s 9586 23933 9642 24733 4 reset
port 12 nsew
rlabel metal4 s 17887 2128 18207 22352 4 VPWR
port 13 nsew
rlabel metal4 s 11110 2128 11430 22352 4 VPWR
port 13 nsew
rlabel metal4 s 4333 2128 4653 22352 4 VPWR
port 13 nsew
rlabel metal5 s 1104 18741 21436 19061 4 VPWR
port 13 nsew
rlabel metal5 s 1104 12032 21436 12352 4 VPWR
port 13 nsew
rlabel metal5 s 1104 5323 21436 5643 4 VPWR
port 13 nsew
rlabel metal4 s 14499 2128 14819 22352 4 VGND
port 14 nsew
rlabel metal4 s 7721 2128 8041 22352 4 VGND
port 14 nsew
rlabel metal5 s 1104 15387 21436 15707 4 VGND
port 14 nsew
rlabel metal5 s 1104 8677 21436 8997 4 VGND
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 22589 24733
<< end >>
