module vm (clk,
    reset,
    VPWR,
    VGND,
    change,
    choice,
    coin,
    out);
 input clk;
 input reset;
 input VPWR;
 input VGND;
 output [1:0] change;
 input [2:0] choice;
 input [1:0] coin;
 output [2:0] out;

 sky130_fd_sc_hd__inv_2 _075_ (.A(reset),
    .Y(_019_));
 sky130_fd_sc_hd__buf_2 _076_ (.A(_019_),
    .X(_020_));
 sky130_fd_sc_hd__buf_2 _077_ (.A(_020_),
    .X(_021_));
 sky130_fd_sc_hd__or2_4 _078_ (.A(coin[0]),
    .B(coin[1]),
    .X(_022_));
 sky130_fd_sc_hd__inv_2 _079_ (.A(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__buf_2 _080_ (.A(\state[7] ),
    .X(_024_));
 sky130_fd_sc_hd__or2_4 _081_ (.A(\state[4] ),
    .B(\state[5] ),
    .X(_025_));
 sky130_fd_sc_hd__or3_4 _082_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(\state[6] ),
    .X(_026_));
 sky130_fd_sc_hd__or4_4 _083_ (.A(_024_),
    .B(_025_),
    .C(\state[2] ),
    .D(_026_),
    .X(_027_));
 sky130_fd_sc_hd__or4_4 _084_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(\state[2] ),
    .D(_025_),
    .X(_028_));
 sky130_fd_sc_hd__or4_4 _085_ (.A(\state[6] ),
    .B(\state[7] ),
    .C(\state[0] ),
    .D(_028_),
    .X(_029_));
 sky130_fd_sc_hd__inv_2 _086_ (.A(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__a21o_4 _087_ (.A1(_023_),
    .A2(_027_),
    .B1(_030_),
    .X(_031_));
 sky130_fd_sc_hd__inv_2 _088_ (.A(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__or2_4 _089_ (.A(change[0]),
    .B(_032_),
    .X(_033_));
 sky130_fd_sc_hd__buf_2 _090_ (.A(coin[0]),
    .X(_034_));
 sky130_fd_sc_hd__inv_2 _091_ (.A(coin[1]),
    .Y(_035_));
 sky130_fd_sc_hd__buf_2 _092_ (.A(_035_),
    .X(_036_));
 sky130_fd_sc_hd__or2_4 _093_ (.A(_034_),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__inv_2 _094_ (.A(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__and2_4 _095_ (.A(coin[0]),
    .B(_035_),
    .X(_039_));
 sky130_fd_sc_hd__inv_2 _096_ (.A(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__or2_4 _097_ (.A(_024_),
    .B(_025_),
    .X(_041_));
 sky130_fd_sc_hd__and3_4 _098_ (.A(_040_),
    .B(_037_),
    .C(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a211o_4 _099_ (.A1(_026_),
    .A2(_038_),
    .B1(_042_),
    .C1(_031_),
    .X(_043_));
 sky130_fd_sc_hd__and3_4 _100_ (.A(_021_),
    .B(_033_),
    .C(_043_),
    .X(_011_));
 sky130_fd_sc_hd__a21oi_4 _101_ (.A1(_036_),
    .A2(_028_),
    .B1(_024_),
    .Y(_044_));
 sky130_fd_sc_hd__or2_4 _102_ (.A(\state[6] ),
    .B(_024_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_4 _103_ (.A1(_045_),
    .A2(_023_),
    .B1(_030_),
    .X(_046_));
 sky130_fd_sc_hd__inv_2 _104_ (.A(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__o21a_4 _105_ (.A1(_039_),
    .A2(_044_),
    .B1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__a21oi_4 _106_ (.A1(_024_),
    .A2(_047_),
    .B1(out[2]),
    .Y(_049_));
 sky130_fd_sc_hd__or3_4 _107_ (.A(reset),
    .B(_048_),
    .C(_049_),
    .X(_050_));
 sky130_fd_sc_hd__inv_2 _108_ (.A(_050_),
    .Y(_010_));
 sky130_fd_sc_hd__a21o_4 _109_ (.A1(_029_),
    .A2(_022_),
    .B1(out[1]),
    .X(_051_));
 sky130_fd_sc_hd__buf_2 _110_ (.A(\state[2] ),
    .X(_052_));
 sky130_fd_sc_hd__and2_4 _111_ (.A(_052_),
    .B(_034_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_4 _112_ (.A1(\state[5] ),
    .A2(_053_),
    .B1(_040_),
    .X(_054_));
 sky130_fd_sc_hd__or3_4 _113_ (.A(\state[1] ),
    .B(_052_),
    .C(\state[4] ),
    .X(_055_));
 sky130_fd_sc_hd__and2_4 _114_ (.A(_023_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__or2_4 _115_ (.A(\state[6] ),
    .B(_046_),
    .X(_057_));
 sky130_fd_sc_hd__or4_4 _116_ (.A(\state[3] ),
    .B(_054_),
    .C(_056_),
    .D(_057_),
    .X(_058_));
 sky130_fd_sc_hd__and3_4 _117_ (.A(_021_),
    .B(_051_),
    .C(_058_),
    .X(_009_));
 sky130_fd_sc_hd__or2_4 _118_ (.A(out[0]),
    .B(_047_),
    .X(_059_));
 sky130_fd_sc_hd__or3_4 _119_ (.A(\state[2] ),
    .B(\state[3] ),
    .C(\state[5] ),
    .X(_060_));
 sky130_fd_sc_hd__and2_4 _120_ (.A(_035_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__o21a_4 _121_ (.A1(\state[4] ),
    .A2(_061_),
    .B1(_040_),
    .X(_062_));
 sky130_fd_sc_hd__o22a_4 _122_ (.A1(\state[1] ),
    .A2(_062_),
    .B1(out[0]),
    .B2(_022_),
    .X(_063_));
 sky130_fd_sc_hd__or2_4 _123_ (.A(_057_),
    .B(_063_),
    .X(_064_));
 sky130_fd_sc_hd__and3_4 _124_ (.A(_021_),
    .B(_059_),
    .C(_064_),
    .X(_008_));
 sky130_fd_sc_hd__inv_2 _125_ (.A(choice[0]),
    .Y(_065_));
 sky130_fd_sc_hd__or3_4 _126_ (.A(choice[2]),
    .B(choice[1]),
    .C(_065_),
    .X(_066_));
 sky130_fd_sc_hd__inv_2 _127_ (.A(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__and3_4 _128_ (.A(_021_),
    .B(\state[0] ),
    .C(_067_),
    .X(_002_));
 sky130_fd_sc_hd__inv_2 _129_ (.A(choice[2]),
    .Y(_068_));
 sky130_fd_sc_hd__and3_4 _130_ (.A(_019_),
    .B(\state[0] ),
    .C(_066_),
    .X(_069_));
 sky130_fd_sc_hd__and4_4 _131_ (.A(_068_),
    .B(choice[1]),
    .C(_069_),
    .D(_065_),
    .X(_001_));
 sky130_fd_sc_hd__and4_4 _132_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(_052_),
    .X(_003_));
 sky130_fd_sc_hd__and4_4 _133_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(\state[4] ),
    .X(_000_));
 sky130_fd_sc_hd__and4_4 _134_ (.A(_068_),
    .B(choice[1]),
    .C(_069_),
    .D(choice[0]),
    .X(_004_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(choice[1]),
    .Y(_070_));
 sky130_fd_sc_hd__and4_4 _136_ (.A(choice[2]),
    .B(_070_),
    .C(_065_),
    .D(_069_),
    .X(_005_));
 sky130_fd_sc_hd__and4_4 _137_ (.A(_034_),
    .B(_036_),
    .C(_020_),
    .D(\state[5] ),
    .X(_071_));
 sky130_fd_sc_hd__and4_4 _138_ (.A(_020_),
    .B(_040_),
    .C(_052_),
    .D(_038_),
    .X(_072_));
 sky130_fd_sc_hd__or2_4 _139_ (.A(_071_),
    .B(_072_),
    .X(_007_));
 sky130_fd_sc_hd__o32a_4 _140_ (.A1(_068_),
    .A2(choice[1]),
    .A3(choice[0]),
    .B1(choice[2]),
    .B2(_070_),
    .X(_073_));
 sky130_fd_sc_hd__or4_4 _141_ (.A(\state[1] ),
    .B(\state[3] ),
    .C(reset),
    .D(_045_),
    .X(_074_));
 sky130_fd_sc_hd__a21oi_4 _142_ (.A1(_052_),
    .A2(_037_),
    .B1(_025_),
    .Y(_013_));
 sky130_fd_sc_hd__or3_4 _143_ (.A(reset),
    .B(_039_),
    .C(_013_),
    .X(_014_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__a211o_4 _145_ (.A1(_069_),
    .A2(_073_),
    .B1(_074_),
    .C1(_015_),
    .X(_006_));
 sky130_fd_sc_hd__or2_4 _146_ (.A(change[1]),
    .B(_032_),
    .X(_016_));
 sky130_fd_sc_hd__and3_4 _147_ (.A(_040_),
    .B(_037_),
    .C(_026_),
    .X(_017_));
 sky130_fd_sc_hd__or2_4 _148_ (.A(_031_),
    .B(_017_),
    .X(_018_));
 sky130_fd_sc_hd__and3_4 _149_ (.A(_021_),
    .B(_016_),
    .C(_018_),
    .X(_012_));
 sky130_fd_sc_hd__dfxtp_4 _150_ (.D(_006_),
    .Q(\state[0] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _151_ (.D(_000_),
    .Q(\state[1] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _152_ (.D(_001_),
    .Q(\state[2] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _153_ (.D(_007_),
    .Q(\state[3] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _154_ (.D(_002_),
    .Q(\state[4] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _155_ (.D(_003_),
    .Q(\state[5] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _156_ (.D(_004_),
    .Q(\state[6] ),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _157_ (.D(_005_),
    .Q(\state[7] ),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _158_ (.D(_008_),
    .Q(out[0]),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _159_ (.D(_009_),
    .Q(out[1]),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _160_ (.D(_010_),
    .Q(out[2]),
    .CLK(clknet_1_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _161_ (.D(_011_),
    .Q(change[0]),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _162_ (.D(_012_),
    .Q(change[1]),
    .CLK(clknet_1_0_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__decap_12 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_23 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_7 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_20 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_82 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_38 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_107 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_77 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_114 ();
endmodule
